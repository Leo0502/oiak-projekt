//: version "2.0.0"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "z80.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 [14:0] w165;    //: /sn:0 {0}(#:-1507,-1232)(-1507,-1203){1}
supply1 w237;    //: /sn:0 {0}(153,-653)(153,-635){1}
//: {2}(151,-633)(135,-633)(135,-606)(142,-606){3}
//: {4}(153,-631)(153,-627){5}
supply1 w132;    //: /sn:0 {0}(-1103,-1290)(-1103,-1315){1}
//: {2}(-1101,-1317)(-1072,-1317)(-1072,-1269)(-1082,-1269){3}
//: {4}(-1103,-1319)(-1103,-1330){5}
supply0 w119;    //: /sn:0 {0}(-1553,-234)(-1553,-211){1}
supply1 w247;    //: /sn:0 {0}(154,-1317)(154,-1303){1}
//: {2}(152,-1301)(138,-1301)(138,-1269)(143,-1269){3}
//: {4}(154,-1299)(154,-1290){5}
supply0 w147;    //: /sn:0 {0}(-1496,-882)(-1509,-882){1}
supply0 w115;    //: /sn:0 {0}(246,-132)(221,-132){1}
supply0 w110;    //: /sn:0 {0}(1509,-66)(1468,-66){1}
supply0 w46;    //: /sn:0 {0}(-1619,-1293)(-1639,-1293){1}
supply1 w263;    //: /sn:0 {0}(153,-1528)(153,-1519){1}
//: {2}(151,-1517)(137,-1517)(137,-1480)(142,-1480){3}
//: {4}(153,-1515)(153,-1501){5}
supply0 w35;    //: /sn:0 {0}(628,-536)(588,-536)(588,-566){1}
//: {2}(590,-568)(628,-568){3}
//: {4}(588,-570)(588,-598){5}
//: {6}(590,-600)(628,-600){7}
//: {8}(588,-602)(588,-630){9}
//: {10}(590,-632)(628,-632){11}
//: {12}(588,-634)(588,-742){13}
//: {14}(590,-744)(628,-744){15}
//: {16}(588,-746)(588,-790){17}
//: {18}(590,-792)(628,-792){19}
//: {20}(588,-794)(588,-968){21}
reg CLR;    //: /sn:0 {0}(-1452,-509)(-1441,-509){1}
supply1 w243;    //: /sn:0 {0}(152,-749)(152,-731){1}
//: {2}(150,-729)(134,-729)(134,-702)(141,-702){3}
//: {4}(152,-727)(152,-723){5}
supply0 w166;    //: /sn:0 {0}(-1488,-1134)(-1504,-1134){1}
reg w92;    //: /sn:0 {0}(261,-182)(271,-182)(271,-142)(221,-142){1}
supply0 w43;    //: /sn:0 {0}(106,-1132)(86,-1132)(86,-1147){1}
supply1 w254;    //: /sn:0 {0}(150,-1422)(150,-1410){1}
//: {2}(148,-1408)(133,-1408)(133,-1374)(139,-1374){3}
//: {4}(150,-1406)(150,-1395){5}
supply1 w26;    //: /sn:0 {0}(153,-1218)(153,-1203){1}
//: {2}(151,-1201)(136,-1201)(136,-1174)(142,-1174){3}
//: {4}(153,-1199)(153,-1195){5}
supply1 w239;    //: /sn:0 {0}(153,-554)(153,-541){1}
//: {2}(151,-539)(138,-539)(138,-512)(142,-512){3}
//: {4}(153,-537)(153,-533){5}
supply1 w241;    //: /sn:0 {0}(153,-465)(153,-450){1}
//: {2}(151,-448)(137,-448)(137,-417)(142,-417){3}
//: {4}(153,-446)(153,-438){5}
supply1 w225;    //: /sn:0 {0}(153,-1029)(153,-1015){1}
//: {2}(151,-1013)(136,-1013)(136,-987)(142,-987){3}
//: {4}(153,-1011)(153,-1008){5}
supply1 w154;    //: /sn:0 {0}(-982,-914)(-990,-914)(-990,-1005){1}
//: {2}(-988,-1007)(-973,-1007){3}
//: {4}(-969,-1007)(-856,-1007){5}
//: {6}(-852,-1007)(-839,-1007){7}
//: {8}(-835,-1007)(-734,-1007){9}
//: {10}(-730,-1007)(-716,-1007){11}
//: {12}(-712,-1007)(-609,-1007){13}
//: {14}(-605,-1007)(-589,-1007){15}
//: {16}(-585,-1007)(-478,-1007){17}
//: {18}(-474,-1007)(-463,-1007){19}
//: {20}(-459,-1007)(-329,-1007){21}
//: {22}(-325,-1007)(-307,-1007)(-307,-841){23}
//: {24}(-327,-1005)(-327,-820)(-318,-820){25}
//: {26}(-461,-1005)(-461,-950){27}
//: {28}(-476,-1005)(-476,-929)(-472,-929){29}
//: {30}(-587,-1005)(-587,-841){31}
//: {32}(-607,-1005)(-607,-820)(-598,-820){33}
//: {34}(-714,-1005)(-714,-935){35}
//: {36}(-732,-1005)(-732,-914)(-725,-914){37}
//: {38}(-837,-1005)(-837,-841){39}
//: {40}(-854,-1005)(-854,-820)(-848,-820){41}
//: {42}(-971,-1005)(-971,-935){43}
//: {44}(-992,-1007)(-1101,-1007){45}
//: {46}(-1105,-1007)(-1126,-1007){47}
//: {48}(-1130,-1007)(-1195,-1007){49}
//: {50}(-1197,-1009)(-1197,-1022){51}
//: {52}(-1197,-1005)(-1197,-841){53}
//: {54}(-1128,-1005)(-1128,-820)(-1114,-820){55}
//: {56}(-1103,-1005)(-1103,-841){57}
supply1 w156;    //: /sn:0 {0}(-1517,-1256)(-1517,-1203){1}
supply1 w131;    //: /sn:0 {0}(-1260,-1290)(-1260,-1313){1}
//: {2}(-1258,-1315)(-1229,-1315)(-1229,-1269)(-1239,-1269){3}
//: {4}(-1260,-1317)(-1260,-1330){5}
supply1 w232;    //: /sn:0 {0}(152,-843)(152,-827){1}
//: {2}(150,-825)(133,-825)(133,-799)(141,-799){3}
//: {4}(152,-823)(152,-820){5}
supply0 w17;    //: /sn:0 {0}(1446,136)(1446,126)(1509,126){1}
//: {2}(1513,126)(1549,126){3}
//: {4}(1511,124)(1511,121)(1525,121){5}
//: {6}(1529,121)(1549,121){7}
//: {8}(1527,119)(1527,62){9}
//: {10}(1527,58)(1527,-14){11}
//: {12}(1525,60)(1522,60)(1522,-14){13}
supply1 w219;    //: /sn:0 {0}(153,-1127)(153,-1113){1}
//: {2}(151,-1111)(135,-1111)(135,-1080)(142,-1080){3}
//: {4}(153,-1109)(153,-1101){5}
supply0 w47;    //: /sn:0 {0}(107,-1434)(82,-1434)(82,-1454){1}
supply1 w146;    //: /sn:0 {0}(-964,-1290)(-964,-1311){1}
//: {2}(-962,-1313)(-933,-1313)(-933,-1269)(-943,-1269){3}
//: {4}(-964,-1315)(-964,-1330){5}
supply0 w160;    //: /sn:0 {0}(1703,-10)(1719,-10){1}
supply1 w231;    //: /sn:0 {0}(153,-937)(153,-921){1}
//: {2}(151,-919)(134,-919)(134,-893)(142,-893){3}
//: {4}(153,-917)(153,-914){5}
wire w16;    //: /sn:0 {0}(1023,-840)(1066,-840){1}
wire w207;    //: /sn:0 {0}(174,-616)(232,-616)(232,-648)(415,-648){1}
//: {2}(419,-648)(522,-648)(522,-648)(628,-648){3}
//: {4}(417,-646)(417,-524)(417,-524)(417,-401){5}
wire w242;    //: /sn:0 {0}(-409,-717)(-409,-401){1}
//: {2}(-407,-399)(42,-399){3}
//: {4}(44,-401)(44,-453){5}
//: {6}(46,-455)(91,-455)(91,-487){7}
//: {8}(44,-457)(44,-652){9}
//: {10}(46,-654)(82,-654)(82,-671){11}
//: {12}(44,-656)(44,-760){13}
//: {14}(46,-762)(76,-762)(76,-777){15}
//: {16}(44,-764)(44,-861){17}
//: {18}(46,-863)(77,-863)(77,-871){19}
//: {20}(44,-865)(44,-1043){21}
//: {22}(46,-1045)(82,-1045)(82,-1057){23}
//: {24}(44,-1047)(44,-1331)(89,-1331)(89,-1348){25}
//: {26}(44,-397)(44,-379)(90,-379)(90,-391){27}
//: {28}(-411,-399)(-527,-399){29}
//: {30}(-529,-401)(-529,-803){31}
//: {32}(-531,-399)(-916,-399){33}
//: {34}(-918,-401)(-918,-729){35}
//: {36}(-920,-399)(-1003,-399)(-1003,-399)(-1073,-399){37}
//: {38}(-1075,-401)(-1075,-551){39}
//: {40}(-1077,-399)(-1151,-399){41}
wire w192;    //: /sn:0 {0}(159,-1258)(159,-1239)(210,-1239){1}
//: {2}(212,-1241)(212,-1344){3}
//: {4}(212,-1348)(212,-1460)(158,-1460)(158,-1469){5}
//: {6}(210,-1346)(155,-1346)(155,-1363){7}
//: {8}(212,-1237)(212,-1151){9}
//: {10}(210,-1149)(158,-1149)(158,-1163){11}
//: {12}(212,-1147)(212,-1060){13}
//: {14}(210,-1058)(158,-1058)(158,-1069){15}
//: {16}(212,-1056)(212,-962){17}
//: {18}(210,-960)(158,-960)(158,-976){19}
//: {20}(212,-958)(212,-865){21}
//: {22}(210,-863)(158,-863)(158,-882){23}
//: {24}(212,-861)(212,-774){25}
//: {26}(210,-772)(157,-772)(157,-788){27}
//: {28}(212,-770)(212,-686){29}
//: {30}(210,-684)(157,-684)(157,-691){31}
//: {32}(212,-682)(212,-580){33}
//: {34}(210,-578)(158,-578)(158,-595){35}
//: {36}(212,-576)(212,-491){37}
//: {38}(210,-489)(158,-489)(158,-501){39}
//: {40}(212,-487)(212,-350)(160,-350){41}
//: {42}(158,-352)(158,-406){43}
//: {44}(156,-350)(-186,-350){45}
//: {46}(-188,-352)(-188,-768)(-300,-768){47}
//: {48}(-302,-770)(-302,-809){49}
//: {50}(-304,-768)(-454,-768){51}
//: {52}(-456,-770)(-456,-918){53}
//: {54}(-458,-768)(-580,-768){55}
//: {56}(-582,-770)(-582,-809){57}
//: {58}(-584,-768)(-707,-768){59}
//: {60}(-709,-770)(-709,-903){61}
//: {62}(-711,-768)(-830,-768){63}
//: {64}(-832,-770)(-832,-809){65}
//: {66}(-834,-768)(-964,-768){67}
//: {68}(-966,-770)(-966,-903){69}
//: {70}(-968,-768)(-1096,-768){71}
//: {72}(-1098,-770)(-1098,-809){73}
//: {74}(-1100,-768)(-1200,-768){75}
//: {76}(-1202,-770)(-1202,-809){77}
//: {78}(-1204,-768)(-1352,-768){79}
//: {80}(-1354,-770)(-1354,-1243)(-1257,-1243){81}
//: {82}(-1253,-1243)(-1100,-1243){83}
//: {84}(-1096,-1243)(-959,-1243)(-959,-1258){85}
//: {86}(-1098,-1245)(-1098,-1258){87}
//: {88}(-1255,-1245)(-1255,-1258){89}
//: {90}(-1356,-768)(-1592,-768){91}
//: {92}(-1594,-770)(-1594,-885){93}
//: {94}(-1592,-887)(-1585,-887){95}
//: {96}(-1596,-887)(-1820,-887)(-1820,-1298)(-1715,-1298){97}
//: {98}(-1594,-766)(-1594,-123)(-1560,-123){99}
//: {100}(-1558,-125)(-1558,-135){101}
//: {102}(-1558,-121)(-1558,-67)(-1613,-67){103}
//: {104}(-188,-348)(-188,-139){105}
//: {106}(-186,-137)(145,-137){107}
//: {108}(-188,-135)(-188,129)(586,129){109}
wire w139;    //: /sn:0 {0}(-890,-1276)(-878,-1276)(-878,-1218)(-1039,-1218){1}
//: {2}(-1041,-1220)(-1041,-1261)(-1016,-1261)(-1016,-1276)(-1026,-1276){3}
//: {4}(-1043,-1218)(-1188,-1218)(-1188,-1276)(-1201,-1276){5}
//: {6}(-1041,-1216)(-1041,-683){7}
wire w58;    //: /sn:0 {0}(163,-438)(163,-447)(195,-447)(195,-543){1}
//: {2}(195,-547)(195,-637){3}
//: {4}(195,-641)(195,-733){5}
//: {6}(195,-737)(195,-825){7}
//: {8}(195,-829)(195,-919){9}
//: {10}(195,-923)(195,-1016){11}
//: {12}(195,-1020)(195,-1112){13}
//: {14}(195,-1116)(195,-1228){15}
//: {16}(195,-1232)(195,-1297){17}
//: {18}(195,-1301)(195,-1403){19}
//: {20}(195,-1407)(195,-1512)(163,-1512)(163,-1501){21}
//: {22}(193,-1405)(160,-1405)(160,-1395){23}
//: {24}(193,-1299)(164,-1299)(164,-1290){25}
//: {26}(193,-1230)(165,-1230){27}
//: {28}(161,-1230)(-67,-1230)(-67,-1048)(-295,-1048){29}
//: {30}(-299,-1048)(-449,-1048){31}
//: {32}(-453,-1048)(-575,-1048){33}
//: {34}(-579,-1048)(-702,-1048){35}
//: {36}(-706,-1048)(-825,-1048){37}
//: {38}(-829,-1048)(-959,-1048){39}
//: {40}(-963,-1048)(-1091,-1048){41}
//: {42}(-1095,-1048)(-1205,-1048){43}
//: {44}(-1209,-1048)(-1370,-1048){45}
//: {46}(-1372,-1050)(-1372,-1301){47}
//: {48}(-1370,-1303)(-1252,-1303){49}
//: {50}(-1248,-1303)(-1095,-1303){51}
//: {52}(-1091,-1303)(-954,-1303)(-954,-1290){53}
//: {54}(-1093,-1301)(-1093,-1290){55}
//: {56}(-1250,-1301)(-1250,-1290){57}
//: {58}(-1374,-1303)(-1639,-1303){59}
//: {60}(-1372,-1046)(-1372,-894){61}
//: {62}(-1374,-892)(-1509,-892){63}
//: {64}(-1372,-890)(-1372,-511){65}
//: {66}(-1374,-509)(-1425,-509){67}
//: {68}(-1372,-507)(-1372,-482)(-1455,-482){69}
//: {70}(-1459,-482)(-1563,-482)(-1563,-211){71}
//: {72}(-1457,-480)(-1457,418)(586,418){73}
//: {74}(-1207,-1046)(-1207,-841){75}
//: {76}(-1093,-1046)(-1093,-841){77}
//: {78}(-961,-1046)(-961,-935){79}
//: {80}(-827,-1046)(-827,-841){81}
//: {82}(-704,-1046)(-704,-935){83}
//: {84}(-577,-1046)(-577,-841){85}
//: {86}(-451,-1046)(-451,-950){87}
//: {88}(-297,-1046)(-297,-841){89}
//: {90}(163,-1228)(163,-1195){91}
//: {92}(193,-1114)(163,-1114)(163,-1101){93}
//: {94}(193,-1018)(163,-1018)(163,-1008){95}
//: {96}(193,-921)(163,-921)(163,-914){97}
//: {98}(193,-827)(162,-827)(162,-820){99}
//: {100}(193,-735)(162,-735)(162,-723){101}
//: {102}(193,-639)(163,-639)(163,-627){103}
//: {104}(193,-545)(163,-545)(163,-533){105}
wire w240;    //: /sn:0 {0}(87,-1057)(87,-1031)(36,-1031){1}
//: {2}(34,-1033)(34,-1239)(93,-1239)(93,-1243){3}
//: {4}(34,-1029)(34,-951){5}
//: {6}(36,-949)(80,-949)(80,-962){7}
//: {8}(34,-947)(34,-566){9}
//: {10}(36,-564)(83,-564)(83,-575){11}
//: {12}(34,-562)(34,-467){13}
//: {14}(36,-465)(86,-465)(86,-487){15}
//: {16}(34,-463)(34,-417){17}
//: {18}(32,-415)(-412,-415){19}
//: {20}(-414,-417)(-414,-717){21}
//: {22}(-416,-415)(-658,-415){23}
//: {24}(-660,-417)(-660,-700){25}
//: {26}(-662,-415)(-911,-415){27}
//: {28}(-913,-417)(-913,-729){29}
//: {30}(-915,-415)(-998,-415)(-998,-415)(-1068,-415){31}
//: {32}(-1070,-417)(-1070,-551){33}
//: {34}(-1072,-415)(-1151,-415){35}
//: {36}(34,-413)(34,-372)(95,-372)(95,-391){37}
wire w88;    //: /sn:0 {0}(-1137,-656)(-1068,-656)(-1068,-572){1}
wire [7:0] w50;    //: /sn:0 {0}(#:1590,224)(1590,234)(1640,234){1}
//: {2}(1642,232)(#:1642,140){3}
//: {4}(1642,236)(1642,515)(182,515)(182,255){5}
//: {6}(184,253)(417,253)(417,253)(#:586,253){7}
//: {8}(182,251)(182,-33){9}
//: {10}(184,-35)(258,-35)(258,46)(#:586,46){11}
//: {12}(182,-37)(182,-91){13}
//: {14}(184,-93)(320,-93)(320,-248)(305,-248){15}
//: {16}(182,-95)(182,-111){17}
//: {18}(182,-115)(#:182,-126){19}
//: {20}(180,-113)(102,-113)(#:102,-171){21}
wire w197;    //: /sn:0 {0}(128,-1279)(143,-1279){1}
wire w81;    //: /sn:0 {0}(-1065,-551)(-1065,-433){1}
//: {2}(-1063,-431)(-1001,-431)(-1001,-431)(-925,-431){3}
//: {4}(-921,-431)(-758,-431)(-758,-857){5}
//: {6}(-923,-433)(-923,-589)(-923,-589)(-923,-729){7}
//: {8}(-1067,-431)(-1151,-431){9}
wire w39;    //: /sn:0 {0}(407,-401)(407,-518){1}
//: {2}(409,-520)(628,-520){3}
//: {4}(405,-520)(243,-520)(243,-427)(174,-427){5}
wire w4;    //: /sn:0 {0}(-1728,-666)(-1821,-666)(-1821,-133)(-1752,-133)(-1752,-156){1}
wire w229;    //: /sn:0 {0}(-800,-878)(-800,-894){1}
//: {2}(-798,-896)(-790,-896){3}
//: {4}(-786,-896)(-631,-896)(-631,-942)(-543,-942){5}
//: {6}(-539,-942)(-517,-942){7}
//: {8}(-541,-944)(-541,-1493)(62,-1493){9}
//: {10}(66,-1493)(96,-1493){11}
//: {12}(64,-1491)(64,-1389){13}
//: {14}(66,-1387)(103,-1387){15}
//: {16}(64,-1385)(64,-1284){17}
//: {18}(66,-1282)(107,-1282){19}
//: {20}(64,-1280)(64,-1189){21}
//: {22}(66,-1187)(102,-1187){23}
//: {24}(64,-1185)(64,-1095){25}
//: {26}(66,-1093)(100,-1093){27}
//: {28}(64,-1091)(64,-1002){29}
//: {30}(66,-1000)(98,-1000){31}
//: {32}(64,-998)(64,-908){33}
//: {34}(66,-906)(95,-906){35}
//: {36}(64,-904)(64,-814){37}
//: {38}(66,-812)(94,-812){39}
//: {40}(64,-810)(64,-717){41}
//: {42}(66,-715)(97,-715){43}
//: {44}(64,-713)(64,-621){45}
//: {46}(66,-619)(98,-619){47}
//: {48}(64,-617)(64,-527){49}
//: {50}(66,-525)(108,-525){51}
//: {52}(64,-523)(64,-430)(106,-430){53}
//: {54}(-788,-894)(-788,-833)(-644,-833){55}
//: {56}(-800,-898)(-800,-927)(-756,-927){57}
wire w56;    //: /sn:0 {0}(-1707,-666)(-1690,-666)(-1690,-802)(-1637,-802){1}
//: {2}(-1633,-802)(-1152,-802)(-1152,-828){3}
//: {4}(-1150,-830)(-1114,-830){5}
//: {6}(-1154,-830)(-1186,-830){7}
//: {8}(-1635,-800)(-1635,-196){9}
wire w123;    //: /sn:0 {0}(1570,124)(1609,124){1}
wire w109;    //: /sn:0 {0}(-1222,-1279)(-1239,-1279){1}
wire w177;    //: /sn:0 {0}(142,-903)(116,-903){1}
wire [7:0] w22;    //: /sn:0 {0}(#:-1528,-1449)(-1528,-1488)(-1529,-1488)(-1529,-1519){1}
//: {2}(#:-1527,-1521)(-1457,-1521)(-1457,-1449){3}
//: {4}(-1531,-1521)(#:-1917,-1521)(-1917,-110)(-1709,-110){5}
//: {6}(-1707,-112)(-1707,-181){7}
//: {8}(-1705,-183)(#:-1651,-183){9}
//: {10}(-1709,-183)(#:-1735,-183){11}
//: {12}(-1707,-108)(-1707,227)(35,227)(#:35,-84){13}
wire [7:0] w3;    //: /sn:0 {0}(#:1177,-667)(1177,-497)(564,-497)(564,170)(#:586,170){1}
wire w128;    //: /sn:0 {0}(-735,-924)(-725,-924){1}
wire w189;    //: /sn:0 {0}(-412,-738)(-412,-828)(-406,-828){1}
wire [7:0] w0;    //: /sn:0 {0}(#:945,129)(985,129)(985,482)(55,482)(55,-84){1}
wire w226;    //: /sn:0 {0}(94,-807)(76,-807)(76,-798){1}
wire w209;    //: /sn:0 {0}(119,-616)(142,-616){1}
wire w20;    //: /sn:0 {0}(-1060,-551)(-1060,-449){1}
//: {2}(-1058,-447)(-1049,-447)(-1049,-447)(-1026,-447){3}
//: {4}(-1022,-447)(-763,-447)(-763,-857){5}
//: {6}(-1024,-449)(-1024,-864){7}
//: {8}(-1062,-447)(-1151,-447){9}
wire w261;    //: /sn:0 {0}(174,-1480)(189,-1480){1}
wire w30;    //: /sn:0 {0}(174,-903)(249,-903)(249,-712)(425,-712){1}
//: {2}(429,-712)(529,-712)(529,-712)(628,-712){3}
//: {4}(427,-710)(427,-412)(427,-412)(427,-401){5}
wire [7:0] w29;    //: /sn:0 {0}(#:1616,-13)(1616,-271)(263,-271){1}
wire w122;    //: /sn:0 {0}(1525,-35)(1525,-53){1}
wire w185;    //: /sn:0 {0}(412,-401)(412,-572)(412,-572)(412,-582){1}
//: {2}(414,-584)(522,-584)(522,-584)(628,-584){3}
//: {4}(410,-584)(240,-584)(240,-522)(174,-522){5}
wire w195;    //: /sn:0 {0}(127,-427)(142,-427){1}
wire [7:0] w42;    //: /sn:0 {0}(#:45,-113)(45,-156)(82,-156)(82,-171){1}
wire w218;    //: /sn:0 {0}(84,-1078)(84,-1088)(100,-1088){1}
wire w152;    //: /sn:0 {0}(-385,-830)(-318,-830){1}
wire w18;    //: /sn:0 {0}(1023,-856)(1066,-856){1}
wire w12;    //: /sn:0 {0}(1023,-808)(1066,-808){1}
wire w19;    //: /sn:0 {0}(209,-303)(-135,-303){1}
//: {2}(-137,-305)(-137,-804)(-435,-804)(-435,-849){3}
//: {4}(-435,-853)(-435,-939)(-440,-939){5}
//: {6}(-437,-851)(-489,-851)(-489,-835)(-484,-835){7}
//: {8}(-137,-301)(-137,-232)(49,-232){9}
wire w178;    //: /sn:0 {0}(173,-799)(188,-799){1}
wire w138;    //: /sn:0 {0}(-1134,-1119)(-1110,-1119)(-1110,-1233)(-1062,-1233)(-1062,-1277){1}
//: {2}(-1060,-1279)(-1047,-1279){3}
//: {4}(-1064,-1279)(-1082,-1279){5}
wire w91;    //: /sn:0 {0}(1023,-760)(1066,-760){1}
wire w180;    //: /sn:0 {0}(-760,-878)(-760,-922)(-756,-922){1}
wire [7:0] w86;    //: /sn:0 {0}(#:1322,-667)(1322,-548){1}
//: {2}(1324,-546)(#:1386,-546){3}
//: {4}(1322,-544)(1322,-474)(1043,-474)(1043,87)(#:945,87){5}
wire [15:0] w31;    //: /sn:0 {0}(#:-1544,-1148)(-1544,-1164)(-1861,-1164)(-1861,-1104){1}
//: {2}(-1859,-1102)(-1548,-1102)(-1548,-1084){3}
//: {4}(-1861,-1100)(-1861,-1040)(-1861,-1040)(-1861,-863){5}
//: {6}(#:-1859,-861)(-1548,-861)(#:-1548,-876){7}
//: {8}(-1861,-859)(-1861,-181)(#:-1770,-181){9}
wire w106;    //: /sn:0 {0}(1739,-482)(1754,-482){1}
wire w104;    //: /sn:0 {0}(1739,-514)(1754,-514){1}
wire w250;    //: /sn:0 {0}(89,-1369)(89,-1382)(103,-1382){1}
wire w116;    //: /sn:0 {0}(1538,-76)(1582,-76)(1582,-43){1}
//: {2}(1584,-41)(1651,-41)(1651,-289){3}
//: {4}(1582,-39)(1582,2)(1592,2){5}
wire [7:0] w32;    //: /sn:0 {0}(#:182,-147)(182,-157){1}
//: {2}(184,-159)(493,-159)(493,-550){3}
//: {4}(#:495,-552)(#:628,-552){5}
//: {6}(493,-554)(493,-614){7}
//: {8}(495,-616)(#:628,-616){9}
//: {10}(#:493,-618)(493,-760)(628,-760){11}
//: {12}(182,-161)(#:182,-216){13}
wire [15:0] w68;    //: /sn:0 {0}(-1593,-1421)(-1533,-1421)(#:-1533,-1443){1}
wire w53;    //: /sn:0 {0}(123,-1184)(142,-1184){1}
wire w8;    //: /sn:0 {0}(1023,-792)(1066,-792){1}
wire [3:0] w140;    //: /sn:0 {0}(1743,-30)(#:1743,-25){1}
wire w230;    //: /sn:0 {0}(108,-520)(88,-520)(88,-508){1}
wire w233;    //: /sn:0 {0}(92,-412)(92,-425)(106,-425){1}
wire w95;    //: /sn:0 {0}(174,-1490)(330,-1490)(330,-888)(628,-888){1}
wire w89;    //: /sn:0 {0}(-1155,-1111)(-1398,-1111)(-1398,-1071)(-1428,-1071){1}
wire [15:0] w44;    //: /sn:0 {0}(#:-1548,-940)(-1548,-897){1}
wire w167;    //: /sn:0 {0}(119,-997)(142,-997){1}
wire [3:0] w67;    //: /sn:0 {0}(1570,50)(#:1570,62)(1727,62)(1727,4){1}
wire w136;    //: /sn:0 {0}(-660,-721)(-660,-828)(-644,-828){1}
wire w134;    //: /sn:0 {0}(-566,-820)(-551,-820){1}
wire w28;    //: /sn:0 {0}(432,-401)(432,-726){1}
//: {2}(434,-728)(628,-728){3}
//: {4}(430,-728)(264,-728)(264,-997)(174,-997){5}
wire w135;    //: /sn:0 {0}(-623,-830)(-598,-830){1}
wire w187;    //: /sn:0 {0}(129,-522)(142,-522){1}
wire [15:0] w14;    //: /sn:0 {0}(#:-1678,-1332)(-1678,-1308){1}
wire [15:0] w45;    //: /sn:0 {0}(#:-1622,-1411)(-1668,-1411)(-1668,-1361){1}
wire w153;    //: /sn:0 {0}(-975,-1269)(-990,-1269){1}
wire [7:0] w41;    //: /sn:0 {0}(#:234,-261)(192,-261)(192,-245){1}
wire w2;    //: /sn:0 {0}(1023,-776)(1066,-776){1}
wire w74;    //: /sn:0 {0}(1023,-712)(1066,-712){1}
wire w120;    //: /sn:0 {0}(56,-187)(69,-187){1}
wire [7:0] w11;    //: /sn:0 {0}(172,-245)(172,-255)(92,-255)(#:92,-200){1}
wire w78;    //: /sn:0 {0}(174,-1080)(189,-1080){1}
wire w155;    //: /sn:0 {0}(-529,-824)(-529,-937)(-517,-937){1}
wire w129;    //: /sn:0 {0}(628,-776)(609,-776)(609,-313)(1654,-313)(1654,-310){1}
wire w105;    //: /sn:0 {0}(1739,-498)(1754,-498){1}
wire w127;    //: /sn:0 {0}(-693,-914)(-678,-914){1}
wire w15;    //: /sn:0 {0}(1023,-824)(1066,-824){1}
wire w55;    //: /sn:0 {0}(-1137,-661)(-1068,-661)(-1068,-820)(-1082,-820){1}
wire w94;    //: /sn:0 {0}(1656,-289)(1656,-280){1}
//: {2}(1654,-278)(600,-278)(600,-872)(628,-872){3}
//: {4}(1656,-276)(1656,2)(1640,2){5}
wire [7:0] w87;    //: /sn:0 {0}(#:1632,16)(1632,80){1}
//: {2}(1632,81)(#:1632,111){3}
wire [15:0] w96;    //: /sn:0 {0}(-1593,-1401)(-1452,-1401)(#:-1452,-1443){1}
wire w76;    //: /sn:0 {0}(70,-229)(159,-229){1}
wire w100;    //: /sn:0 {0}(1023,-888)(1066,-888){1}
wire w99;    //: /sn:0 {0}(1023,-872)(1066,-872){1}
wire w125;    //: /sn:0 {0}(230,-300)(247,-300)(247,-284){1}
wire w40;    //: /sn:0 {0}(174,-1174)(189,-1174){1}
wire [15:0] w13;    //: /sn:0 {0}(#:-1688,-1361)(-1688,-1376)(-1734,-1376){1}
//: {2}(-1736,-1378)(-1736,-1491)(-1539,-1491){3}
//: {4}(-1538,-1491)(-1448,-1491){5}
//: {6}(-1447,-1491)(-1342,-1491){7}
//: {8}(-1736,-1374)(-1736,-1264)(-1680,-1264){9}
//: {10}(-1678,-1266)(#:-1678,-1287){11}
//: {12}(-1678,-1262)(-1678,-999)(-1558,-999)(-1558,-969){13}
wire w6;    //: /sn:0 {0}(628,-824)(288,-824)(288,-1184)(174,-1184){1}
wire w7;    //: /sn:0 {0}(516,87)(586,87){1}
wire [2:0] w143;    //: /sn:0 {0}(#:586,294)(-511,294)(-511,294)(-1672,294){1}
wire w65;    //: /sn:0 {0}(-803,-857)(-803,-847)(-818,-847)(-818,-924)(-936,-924){1}
//: {2}(-940,-924)(-950,-924){3}
//: {4}(-938,-922)(-938,-778)(-175,-778)(-175,-186){5}
//: {6}(-173,-184)(35,-184){7}
//: {8}(-175,-182)(-175,-98)(-20,-98){9}
wire w34;    //: /sn:0 {0}(1767,-10)(1777,-10)(1777,-395)(618,-395)(618,-680)(628,-680){1}
wire w175;    //: /sn:0 {0}(-918,-750)(-918,-828)(-912,-828){1}
wire w59;    //: /sn:0 {0}(-1020,-927)(-1065,-927){1}
//: {2}(-1067,-929)(-1067,-1205)(-868,-1205)(-868,-1281)(-890,-1281){3}
//: {4}(-1067,-925)(-1067,-835){5}
//: {6}(-1065,-833)(-912,-833){7}
//: {8}(-1067,-831)(-1067,-830)(-1082,-830){9}
wire [15:0] w158;    //: /sn:0 {0}(#:-1528,-1119)(-1528,-1084){1}
wire w252;    //: /sn:0 {0}(171,-1374)(186,-1374){1}
wire [2:0] w25;    //: /sn:0 {0}(-1672,377)(-511,377)(-511,377)(#:586,377){1}
wire w72;    //: /sn:0 {0}(-463,-832)(-444,-832)(-444,-833)(-406,-833){1}
wire w186;    //: /sn:0 {0}(174,-512)(189,-512){1}
wire w176;    //: /sn:0 {0}(174,-893)(189,-893){1}
wire w142;    //: /sn:0 {0}(-472,-939)(-496,-939){1}
wire w36;    //: /sn:0 {0}(173,-809)(236,-809)(236,-696)(628,-696){1}
wire [7:0] w82;    //: /sn:0 {0}(#:-1447,-1487)(-1447,-1449){1}
wire w60;    //: /sn:0 {0}(35,-189)(-159,-189){1}
//: {2}(-161,-191)(-161,-787)(-796,-787){3}
//: {4}(-798,-789)(-798,-828){5}
//: {6}(-798,-832)(-798,-857){7}
//: {8}(-800,-830)(-816,-830){9}
//: {10}(-800,-787)(-1681,-787)(-1681,-661)(-1707,-661){11}
//: {12}(-161,-187)(-161,-103)(-20,-103){13}
wire w124;    //: /sn:0 {0}(1,-100)(22,-100){1}
wire w148;    //: /sn:0 {0}(-286,-820)(-271,-820){1}
wire w71;    //: /sn:0 {0}(-1271,-1269)(-1286,-1269){1}
wire [7:0] w112;    //: /sn:0 {0}(#:1590,175)(1590,150)(1622,150)(1622,140){1}
wire w210;    //: /sn:0 {0}(118,-712)(141,-712){1}
wire w235;    //: /sn:0 {0}(82,-692)(82,-710)(97,-710){1}
wire w141;    //: /sn:0 {0}(-440,-929)(-425,-929){1}
wire w227;    //: /sn:0 {0}(83,-596)(83,-614)(98,-614){1}
wire w37;    //: /sn:0 {0}(537,335)(-685,335)(-685,-922){1}
//: {2}(-685,-926)(-685,-1104)(-1078,-1104){3}
//: {4}(-1082,-1104)(-1123,-1104)(-1123,-1104)(-1134,-1104){5}
//: {6}(-1080,-1102)(-1080,-1072)(-1275,-1072){7}
//: {8}(-687,-924)(-693,-924){9}
wire w214;    //: /sn:0 {0}(173,-702)(188,-702){1}
wire [15:0] w168;    //: /sn:0 {0}(#:-1512,-1197)(-1512,-1148){1}
wire w66;    //: /sn:0 {0}(-950,-914)(-935,-914){1}
wire w73;    //: /sn:0 {0}(558,335)(586,335){1}
wire w10;    //: /sn:0 {0}(628,-808)(439,-808){1}
//: {2}(435,-808)(276,-808)(276,-1090)(174,-1090){3}
//: {4}(437,-806)(437,-401){5}
wire [7:0] w23;    //: /sn:0 {0}(#:-1538,-1487)(-1538,-1449){1}
wire w63;    //: /sn:0 {0}(-1275,-1082)(-1265,-1082)(-1265,-1095)(-1297,-1095)(-1297,-1277){1}
//: {2}(-1295,-1279)(-1271,-1279){3}
//: {4}(-1299,-1279)(-1462,-1279)(-1462,-953)(-1525,-953){5}
wire w211;    //: /sn:0 {0}(124,-1384)(139,-1384){1}
wire w179;    //: /sn:0 {0}(141,-809)(115,-809){1}
wire w70;    //: /sn:0 {0}(-1024,-885)(-1024,-922)(-1020,-922){1}
wire w111;    //: /sn:0 {0}(427,-346)(427,-380){1}
wire [7:0] w84;    //: /sn:0 {0}(#:284,-251)(263,-251){1}
wire w24;    //: /sn:0 {0}(628,-840)(444,-840){1}
//: {2}(440,-840)(303,-840)(303,-1279)(175,-1279){3}
//: {4}(442,-838)(442,-401){5}
wire w130;    //: /sn:0 {0}(-1570,-1366)(-1551,-1366)(-1551,-1344){1}
//: {2}(-1549,-1342)(-1144,-1342)(-1144,-1281){3}
//: {4}(-1142,-1279)(-1114,-1279){5}
//: {6}(-1146,-1279)(-1156,-1279)(-1156,-1281)(-1201,-1281){7}
//: {8}(-1553,-1342)(-1568,-1342){9}
wire [15:0] w21;    //: /sn:0 {0}(#:-1538,-1055)(-1538,-969){1}
wire w1;    //: /sn:0 {0}(-1332,-926)(-1332,-1074)(-1313,-1074){1}
//: {2}(-1309,-1074)(-1296,-1074){3}
//: {4}(-1311,-1072)(-1311,-830)(-1218,-830){5}
wire w121;    //: /sn:0 {0}(209,-298)(-147,-298){1}
//: {2}(-149,-300)(-149,-796)(-499,-796)(-499,-828){3}
//: {4}(-497,-830)(-484,-830){5}
//: {6}(-501,-830)(-566,-830){7}
//: {8}(-149,-296)(-149,-227)(49,-227){9}
wire w194;    //: /sn:0 {0}(174,-417)(189,-417){1}
wire w246;    //: /sn:0 {0}(93,-1264)(93,-1277)(107,-1277){1}
wire w224;    //: /sn:0 {0}(95,-901)(77,-901)(77,-892){1}
wire w200;    //: /sn:0 {0}(175,-1269)(190,-1269){1}
wire w182;    //: /sn:0 {0}(-1552,-1134)(-1567,-1134){1}
wire [7:0] w144;    //: /sn:0 {0}(#:-1548,-173)(-1508,-173){1}
//: {2}(-1504,-173)(-1432,-173)(-1432,-447)(#:-1400,-447){3}
//: {4}(-1506,-171)(-1506,-112)(-1674,-112){5}
//: {6}(-1676,-114)(-1676,-163)(-1651,-163){7}
//: {8}(-1676,-110)(-1676,293){9}
//: {10}(-1676,294)(-1676,376){11}
//: {12}(-1676,377)(-1676,397){13}
wire w98;    //: /sn:0 {0}(-1158,-659)(-1266,-659)(-1266,-1067)(-1275,-1067){1}
wire w103;    //: /sn:0 {0}(1739,-530)(1754,-530){1}
wire w52;    //: /sn:0 {0}(-1332,-910)(-1332,-820)(-1218,-820){1}
wire w27;    //: /sn:0 {0}(586,211)(427,211)(427,-325)(-71,-325)(-71,-815)(-119,-815){1}
//: {2}(-121,-817)(-121,-830)(-228,-830){3}
//: {4}(-230,-832)(-230,-1109)(-1093,-1109){5}
//: {6}(-1097,-1109)(-1130,-1109)(-1130,-1109)(-1134,-1109){7}
//: {8}(-1095,-1107)(-1095,-1077)(-1275,-1077){9}
//: {10}(-232,-830)(-286,-830){11}
//: {12}(-121,-813)(-121,87)(495,87){13}
wire w150;    //: /sn:0 {0}(-891,-830)(-881,-830){1}
//: {2}(-877,-830)(-848,-830){3}
//: {4}(-879,-828)(-879,-794)(-1397,-794)(-1397,-1066)(-1428,-1066){5}
wire w113;    //: /sn:0 {0}(-816,-820)(-801,-820){1}
wire w215;    //: /sn:0 {0}(86,-1168)(86,-1182)(102,-1182){1}
wire w118;    //: /sn:0 {0}(174,-987)(189,-987){1}
wire [7:0] w33;    //: /sn:0 {0}(#:1600,16)(1600,46)(1570,46){1}
//: {2}(1569,46)(965,46){3}
//: {4}(963,44)(963,-253)(305,-253){5}
//: {6}(961,46)(#:945,46){7}
wire w163;    //: /sn:0 {0}(-1449,-1068)(-1515,-1068){1}
wire w69;    //: /sn:0 {0}(-999,-924)(-982,-924){1}
wire [7:0] w145;    //: /sn:0 {0}(-1569,-173)(#:-1622,-173){1}
wire w48;    //: /sn:0 {0}(-1151,-367)(-1129,-367)(-1129,-343){1}
wire w257;    //: /sn:0 {0}(82,-1475)(82,-1488)(96,-1488){1}
wire w149;    //: /sn:0 {0}(-1591,-1369)(-1609,-1369)(-1609,-1388){1}
wire w126;    //: /sn:0 {0}(-1186,-820)(-1170,-820){1}
wire w90;    //: /sn:0 {0}(1023,-744)(1066,-744){1}
wire w85;    //: /sn:0 {0}(1023,-728)(1066,-728){1}
wire [3:0] w61;    //: /sn:0 {0}(#:1636,81)(1759,81)(1759,4){1}
wire w5;    //: /sn:0 {0}(117,-1490)(142,-1490){1}
wire w137;    //: /sn:0 {0}(-1114,-1269)(-1129,-1269){1}
wire w38;    //: /sn:0 {0}(-1041,-662)(-1041,-383)(-1151,-383){1}
wire w102;    //: /sn:0 {0}(1509,-86)(1499,-86)(1499,-436)(1762,-436)(1762,-546)(1739,-546){1}
wire w64;    //: /sn:0 {0}(-1707,-671)(-1698,-671)(-1698,-951)(-1594,-951)(-1594,-1343){1}
//: {2}(-1592,-1345)(-1589,-1345){3}
//: {4}(-1596,-1345)(-1655,-1345){5}
wire w9;    //: /sn:0 {0}(422,-401)(422,-662){1}
//: {2}(424,-664)(628,-664){3}
//: {4}(420,-664)(226,-664)(226,-712)(173,-712){5}
wire w221;    //: /sn:0 {0}(80,-983)(80,-995)(98,-995){1}
wire w208;    //: /sn:0 {0}(174,-606)(189,-606){1}
wire w107;    //: /sn:0 {0}(1739,-466)(1754,-466){1}
wire w133;    //: /sn:0 {0}(-1568,-1347)(-1546,-1347){1}
//: {2}(-1542,-1347)(-990,-1347)(-990,-1281){3}
//: {4}(-988,-1279)(-975,-1279){5}
//: {6}(-992,-1279)(-999,-1279)(-999,-1281)(-1026,-1281){7}
//: {8}(-1544,-1349)(-1544,-1371)(-1570,-1371){9}
wire w93;    //: /sn:0 {0}(171,-1384)(316,-1384)(316,-856)(445,-856){1}
//: {2}(449,-856)(628,-856){3}
//: {4}(447,-854)(447,-401){5}
wire w157;    //: /sn:0 {0}(-1134,-1114)(-1102,-1114)(-1102,-1226)(-921,-1226)(-921,-1277){1}
//: {2}(-919,-1279)(-911,-1279){3}
//: {4}(-923,-1279)(-943,-1279){5}
wire w79;    //: /sn:0 {0}(121,-1090)(142,-1090){1}
//: enddecls

  //: joint g8 (w56) @(-1635, -802) /w:[ 2 -1 1 8 ]
  //: joint g164 (w192) @(-456, -768) /w:[ 51 52 54 -1 ]
  //: joint g312 (w192) @(212, -863) /w:[ -1 21 22 24 ]
  _GGJKFF #(10, 10, 20) r_DB (.Q(w65), ._Q(w66), .J(w69), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-966,-919) /w:[ 3 0 1 0 43 79 69 ] /mi:0
  //: joint g224 (w157) @(-921, -1279) /w:[ 2 -1 4 1 ]
  _GGJKFF #(10, 10, 20) DB_r (.Q(w37), ._Q(w127), .J(w128), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-709,-919) /w:[ 9 0 1 37 35 83 61 ] /mi:0
  //: joint g258 (w219) @(153, -1111) /w:[ -1 1 2 4 ]
  _GGJKFF #(10, 10, 20) x1_in_01 (.Q(w6), ._Q(w40), .J(w53), .K(w26), .PRE(w26), .CLR(w58), .CK(w192));   //: @(158,-1179) /w:[ 1 0 1 3 5 91 11 ] /mi:0
  //: joint g226 (w139) @(-1041, -1218) /w:[ 1 2 4 6 ]
  //: joint g243 (w26) @(153, -1201) /w:[ -1 1 2 4 ]
  //: VDD g92 (w219) @(164,-1127) /sn:0 /w:[ 0 ]
  _GGXOR2 #(8) g198 (.I0(w116), .I1(w94), .Z(w129));   //: @(1654,-300) /sn:0 /R:1 /w:[ 3 0 1 ]
  //: VDD g30 (w154) @(-1186,-1022) /sn:0 /w:[ 51 ]
  //: joint g74 (w263) @(153, -1517) /w:[ -1 1 2 4 ]
  //: joint g130 (w27) @(-230, -830) /w:[ 3 4 10 -1 ]
  //: joint g1 (w58) @(-1372, -892) /w:[ -1 61 62 64 ]
  //: joint g183 (w19) @(-137, -303) /w:[ 1 2 -1 8 ]
  _GGREG16 #(10, 10, 20) PC (.Q(w31), .D(w44), .EN(w147), .CLR(w58), .CK(w192));   //: @(-1548,-887) /w:[ 7 1 1 63 95 ]
  //: joint g111 (w154) @(-732, -1007) /w:[ 10 -1 9 36 ]
  //: VDD g253 (w254) @(161,-1422) /sn:0 /w:[ 0 ]
  _GGJKFF #(10, 10, 20) x6_set_b (.Q(w185), ._Q(w186), .J(w187), .K(w239), .PRE(w239), .CLR(w58), .CK(w192));   //: @(158,-517) /w:[ 5 0 1 3 5 105 39 ] /mi:0
  //: joint g260 (w242) @(-409, -399) /w:[ 2 1 28 -1 ]
  _GGAND2 #(6) g274 (.I0(w229), .I1(w226), .Z(w179));   //: @(105,-809) /sn:0 /w:[ 39 0 1 ]
  _GGOR2 #(6) g179 (.I0(w19), .I1(w121), .Z(w76));   //: @(60,-229) /sn:0 /w:[ 9 9 0 ]
  _GGAND2 #(6) g70 (.I0(w229), .I1(w224), .Z(w177));   //: @(106,-903) /sn:0 /w:[ 35 0 1 ]
  //: VDD g206 (w132) @(-1092,-1330) /sn:0 /w:[ 5 ]
  //: joint g149 (w154) @(-837, -1007) /w:[ 8 -1 7 38 ]
  //: GROUND g10 (w115) @(252,-132) /sn:0 /R:1 /w:[ 0 ]
  _GGOR3 #(8) g25 (.I0(w81), .I1(w242), .I2(w240), .Z(w175));   //: @(-918,-740) /sn:0 /R:1 /w:[ 7 35 29 0 ]
  //: joint g220 (w130) @(-1144, -1279) /w:[ 4 3 6 -1 ]
  _GGMUX2x8 #(8, 8) g64 (.I0(w50), .I1(w42), .S(w120), .Z(w11));   //: @(92,-187) /sn:0 /R:2 /w:[ 21 1 1 1 ] /ss:1 /do:0
  //: VDD g49 (w156) @(-1506,-1256) /sn:0 /w:[ 0 ]
  _GGJKFF #(10, 10, 20) AND_DB_DB (.Q(w19), ._Q(w141), .J(w142), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-456,-934) /w:[ 5 0 0 29 27 87 53 ] /mi:0
  //: joint g270 (w229) @(64, -525) /w:[ 50 49 -1 52 ]
  //: joint g35 (w58) @(-577, -1048) /w:[ 33 -1 34 84 ]
  _GGAND2 #(6) g181 (.I0(w19), .I1(!w121), .Z(w125));   //: @(220,-300) /sn:0 /w:[ 0 0 0 ]
  //: joint g192 (w50) @(182, 253) /w:[ 6 8 -1 5 ]
  //: joint g67 (w192) @(-302, -768) /w:[ 47 48 50 -1 ]
  //: GROUND g85 (w166) @(-1482,-1134) /sn:0 /R:1 /w:[ 0 ]
  //: joint g126 (w81) @(-1065, -431) /w:[ 2 1 8 -1 ]
  //: LED g234 (w140) @(1743,-37) /sn:0 /w:[ 0 ] /type:1
  //: joint g33 (w154) @(-971, -1007) /w:[ 4 -1 3 42 ]
  //: joint g54 (w94) @(1656, -278) /w:[ -1 1 2 4 ]
  //: joint g300 (w185) @(412, -584) /w:[ 2 -1 4 1 ]
  _GGAND2 #(4) g132 (.I0(!w88), .I1(!w55), .Z(w98));   //: @(-1148,-659) /sn:0 /R:2 /w:[ 0 0 0 ]
  //: joint g163 (w192) @(-582, -768) /w:[ 55 56 58 -1 ]
  _GGOR1 #(1) g222 (.I0(w38), .Z(w139));   //: @(-1041,-673) /sn:0 /R:1 /w:[ 0 7 ]
  _GGAND2 #(6) g217 (.I0(w139), .I1(w130), .Z(w109));   //: @(-1212,-1279) /sn:0 /R:2 /w:[ 5 7 0 ]
  //: joint g12 (w144) @(-1506, -173) /w:[ 2 -1 1 4 ]
  //: joint g106 (w58) @(163, -1230) /w:[ 27 -1 28 90 ]
  //: joint g298 (w9) @(422, -664) /w:[ 2 -1 4 1 ]
  _GGADD4 #(36, 38, 30, 32) g230 (.A(w61), .B(w67), .S(w140), .CI(w160), .CO(w34));   //: @(1743,-12) /sn:0 /R:2 /w:[ 1 1 1 1 0 ]
  //: joint g194 (w50) @(182, -113) /w:[ -1 18 20 17 ]
  //: joint g177 (w121) @(-499, -830) /w:[ 4 -1 6 3 ]
  //: joint g307 (w192) @(212, -1239) /w:[ -1 2 1 8 ]
  //: joint g228 (w116) @(1582, -41) /w:[ 2 1 -1 4 ]
  //: frame g196 @(279,-290) /sn:0 /wi:56 /ht:68 /tx:"AND"
  //: joint g19 (w81) @(-923, -431) /w:[ 4 6 3 -1 ]
  _GGAND2 #(6) g114 (.I0(w59), .I1(w70), .Z(w69));   //: @(-1009,-924) /sn:0 /w:[ 0 1 0 ]
  _GGJKFF #(10, 10, 20) x0_set_b (.Q(w24), ._Q(w200), .J(w197), .K(w247), .PRE(w247), .CLR(w58), .CK(w192));   //: @(159,-1274) /w:[ 3 0 1 3 5 25 0 ] /mi:0
  _GGOR4 #(10) g125 (.I0(w98), .I1(w37), .I2(w27), .I3(w63), .Z(w1));   //: @(-1286,-1074) /sn:0 /R:2 /w:[ 1 7 9 0 3 ]
  //: joint g281 (w242) @(44, -399) /w:[ -1 4 3 26 ]
  //: VDD g93 (w225) @(164,-1029) /sn:0 /w:[ 0 ]
  _GGJKFF #(10, 10, 20) ADDR_BUS_PC (.Q(w63), ._Q(w71), .J(w109), .K(w131), .PRE(w131), .CLR(w58), .CK(w192));   //: @(-1255,-1274) /w:[ 3 0 1 3 0 57 89 ] /mi:1
  //: GROUND g63 (w165) @(-1507,-1238) /sn:0 /R:2 /w:[ 0 ]
  //: joint g100 (w247) @(154, -1301) /w:[ -1 1 2 4 ]
  //: joint g215 (w133) @(-1544, -1347) /w:[ 2 8 1 -1 ]
  _GGOR2 #(6) g211 (.I0(w130), .I1(w133), .Z(w64));   //: @(-1579,-1345) /sn:0 /R:2 /w:[ 9 0 3 ]
  //: joint g0 (w150) @(-879, -830) /w:[ 2 -1 1 4 ]
  //: joint g101 (w35) @(588, -744) /w:[ 14 16 -1 13 ]
  //: joint g244 (w58) @(195, -545) /w:[ -1 2 104 1 ]
  //: joint g262 (w237) @(153, -633) /w:[ -1 1 2 4 ]
  _GGJKFF #(10, 10, 20) addr_1_half (.Q(w133), ._Q(w153), .J(w157), .K(w146), .PRE(w146), .CLR(w58), .CK(w192));   //: @(-959,-1274) /w:[ 5 0 5 3 0 53 85 ] /mi:1
  registers g37 (.Accumulator_input(w50), .Accumulator_input_choose(w7), .Clock(w192), .Flag_input(w3), .Flag_input_choose(w27), .Register_input(w50), .Register_input_choose(w143), .Register_input_dec(w73), .Register_output_choose1(w25), ._CLR(w58), .Accumulator_output(w33), .Flag_output(w86), .Register_output1(w0));   //: @(587, 5) /sz:(357, 455) /sn:0 /p:[ Li0>11 Li1>1 Li2>109 Li3>1 Li4>0 Li5>7 Li6>0 Li7>1 Li8>1 Li9>73 Ro0<7 Ro1<5 Ro2<0 ]
  _GGOR1 #(1) g120 (.I0(w37), .Z(w73));   //: @(548,335) /sn:0 /w:[ 0 0 ]
  _GGOR2 #(6) g76 (.I0(w242), .I1(w240), .Z(w218));   //: @(84,-1068) /sn:0 /R:1 /w:[ 23 0 0 ]
  _GGJKFF #(10, 10, 20) read_OP (.Q(w56), ._Q(w126), .J(w1), .K(w52), .PRE(w58), .CLR(w154), .CK(w192));   //: @(-1202,-825) /w:[ 7 0 5 1 75 53 77 ] /mi:0
  _GGOR1 #(1) g75 (.I0(w43), .Z(w215));   //: @(86,-1158) /sn:0 /R:1 /w:[ 1 0 ]
  //: GROUND g152 (w147) @(-1490,-882) /sn:0 /R:1 /w:[ 0 ]
  //: joint g267 (w58) @(195, -1299) /w:[ -1 18 24 17 ]
  //: joint g44 (w229) @(64, -1387) /w:[ 14 13 -1 16 ]
  //: frame g159 @(-1844,-230) /sn:0 /wi:120 /ht:108 /tx:""
  //: joint g3 (w58) @(-1457, -482) /w:[ 69 -1 70 72 ]
  //: joint g16 (w17) @(1527, 60) /w:[ -1 10 12 9 ]
  //: joint g47 (w229) @(64, -1493) /w:[ 10 -1 9 12 ]
  //: joint g143 (w56) @(-1152, -830) /w:[ 4 -1 6 3 ]
  _GGOR2 #(6) g26 (.I0(w20), .I1(w81), .Z(w180));   //: @(-760,-868) /sn:0 /R:1 /w:[ 5 5 0 ]
  //: joint g109 (w154) @(-476, -1007) /w:[ 18 -1 17 28 ]
  //: joint g284 (w242) @(44, -455) /w:[ 6 8 -1 5 ]
  //: joint g302 (w192) @(-188, -350) /w:[ 45 46 -1 104 ]
  //: joint g158 (w60) @(-798, -787) /w:[ 3 4 10 -1 ]
  _GGNBUF #(2) g23 (.I(w1), .Z(w52));   //: @(-1332,-920) /sn:0 /R:3 /w:[ 0 0 ]
  //: joint g309 (w192) @(212, -1149) /w:[ -1 9 10 12 ]
  //: joint g86 (w192) @(-1098, -768) /w:[ 71 72 74 -1 ]
  _GGOR1 #(1) g127 (.I0(w27), .Z(w7));   //: @(506,87) /sn:0 /w:[ 13 0 ]
  //: joint g39 (w242) @(-1075, -399) /w:[ 37 38 40 -1 ]
  //: joint g104 (w242) @(-918, -399) /w:[ 33 34 36 -1 ]
  //: joint g24 (w20) @(-1024, -447) /w:[ 4 6 3 -1 ]
  //: LED g316 (w48) @(-1129,-336) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: joint g310 (w192) @(212, -1058) /w:[ -1 13 14 16 ]
  //: joint g121 (w59) @(-1067, -833) /w:[ 6 5 -1 8 ]
  //: joint g110 (w154) @(-607, -1007) /w:[ 14 -1 13 32 ]
  _GGAND2 #(6) g60 (.I0(w229), .I1(w221), .Z(w167));   //: @(109,-997) /sn:0 /w:[ 31 1 0 ]
  _GGAND2 #(6) g250 (.I0(w229), .I1(w250), .Z(w211));   //: @(114,-1384) /sn:0 /w:[ 15 1 0 ]
  //: joint g289 (w240) @(34, -564) /w:[ 10 9 -1 12 ]
  _GGJKFF #(10, 10, 20) DB_A (.Q(w27), ._Q(w148), .J(w152), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-302,-825) /w:[ 11 0 1 25 23 89 49 ] /mi:0
  _GGOR2 #(6) g82 (.I0(w60), .I1(w65), .Z(w120));   //: @(46,-187) /sn:0 /w:[ 0 7 0 ]
  _GGOR1 #(1) g248 (.I0(w240), .Z(w246));   //: @(93,-1254) /sn:0 /R:1 /w:[ 3 0 ]
  //: VDD g257 (w263) @(164,-1528) /sn:0 /w:[ 0 ]
  _GGJKFF #(10, 10, 20) x2_set_par (.Q(w30), ._Q(w176), .J(w177), .K(w231), .PRE(w231), .CLR(w58), .CK(w192));   //: @(158,-898) /w:[ 0 0 0 3 5 97 23 ] /mi:0
  //: joint g306 (w192) @(212, -684) /w:[ -1 29 30 32 ]
  //: joint g272 (w229) @(64, -715) /w:[ 42 41 -1 44 ]
  //: VDD g94 (w231) @(164,-937) /sn:0 /w:[ 0 ]
  //: joint g245 (w58) @(195, -639) /w:[ -1 4 102 3 ]
  _GGMUX2x8 #(8, 8) g107 (.I0(w0), .I1(w22), .S(w124), .Z(w42));   //: @(45,-100) /sn:0 /R:2 /w:[ 1 13 1 0 ] /ss:1 /do:0
  assign w68 = {w22, w23}; //: CONCAT g166  @(-1533,-1444) /sn:0 /R:3 /w:[ 1 0 1 ] /dr:0 /tp:0 /drp:1
  //: joint g216 (w13) @(-1678, -1264) /w:[ -1 10 9 12 ]
  //: joint g301 (w39) @(407, -520) /w:[ 2 -1 4 1 ]
  assign w168 = {w165, w156}; //: CONCAT g68  @(-1512,-1198) /sn:0 /R:3 /w:[ 0 1 1 ] /dr:0 /tp:0 /drp:1
  //: joint g133 (w240) @(-660, -415) /w:[ 23 24 26 -1 ]
  //: joint g263 (w239) @(153, -539) /w:[ -1 1 2 4 ]
  _GGNBUF #(2) g22 (.I(CLR), .Z(w58));   //: @(-1435,-509) /sn:0 /w:[ 1 67 ]
  //: joint g31 (w154) @(-990, -1007) /w:[ 2 -1 44 1 ]
  //: joint g225 (w59) @(-1067, -927) /w:[ 1 2 -1 4 ]
  _GGJKFF #(10, 10, 20) x4_in_01 (.Q(w36), ._Q(w178), .J(w179), .K(w232), .PRE(w232), .CLR(w58), .CK(w192));   //: @(157,-804) /w:[ 0 0 0 3 5 99 27 ] /mi:0
  //: joint g87 (w32) @(493, -616) /w:[ 8 10 -1 7 ]
  //: GROUND g231 (w160) @(1697,-10) /sn:0 /R:3 /w:[ 0 ]
  //: joint g283 (w240) @(34, -465) /w:[ 14 13 -1 16 ]
  //: joint g317 (w64) @(-1594, -1345) /w:[ 2 -1 4 1 ]
  //: joint g83 (w254) @(150, -1408) /w:[ -1 1 2 4 ]
  _GGMUX2x16 #(8, 8) g41 (.I0(w31), .I1(w158), .S(w163), .Z(w21));   //: @(-1538,-1068) /sn:0 /w:[ 3 1 1 0 ] /ss:1 /do:0
  //: joint g203 (w58) @(-1250, -1303) /w:[ 50 -1 49 56 ]
  //: joint g42 (w31) @(-1861, -861) /w:[ 6 5 -1 8 ]
  //: joint g138 (w192) @(-1202, -768) /w:[ 75 76 78 -1 ]
  _GGAND2 #(6) g213 (.I0(!w130), .I1(w133), .Z(w149));   //: @(-1581,-1369) /sn:0 /R:2 /w:[ 0 9 0 ]
  //: joint g264 (w241) @(153, -448) /w:[ -1 1 2 4 ]
  //: joint g293 (w24) @(442, -840) /w:[ 1 -1 2 4 ]
  _GGJKFF #(10, 10, 20) x0_in_01 (.Q(w95), ._Q(w261), .J(w5), .K(w263), .PRE(w263), .CLR(w58), .CK(w192));   //: @(158,-1485) /w:[ 0 0 1 3 5 21 5 ] /mi:0
  assign w96 = {w82, w22}; //: CONCAT g167  @(-1452,-1444) /sn:0 /R:3 /w:[ 1 1 3 ] /dr:0 /tp:0 /drp:1
  //: joint g66 (w240) @(-1070, -415) /w:[ 31 32 34 -1 ]
  //: GROUND g151 (w119) @(-1553,-240) /sn:0 /R:2 /w:[ 0 ]
  _GGMUX2x16 #(8, 8) g153 (.I0(w21), .I1(w13), .S(w63), .Z(w44));   //: @(-1548,-953) /sn:0 /w:[ 1 13 5 0 ] /ss:1 /do:1
  //: joint g146 (w154) @(-461, -1007) /w:[ 20 -1 19 26 ]
  //: joint g162 (w192) @(-709, -768) /w:[ 59 60 62 -1 ]
  //: joint g318 (w27) @(-121, -815) /w:[ 1 2 -1 12 ]
  flags_status g46 (.flags_in(w86), .Flag_7_sign(w107), .Flag_6_zero(w106), .Flag_4_halfcarry(w105), .Flag_2_parity_overflow(w104), .Flag_1_substract(w103), .Flag_0_carry(w102));   //: @(1387, -562) /sz:(351, 112) /sn:0 /p:[ Li0>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 ]
  //: joint g34 (w58) @(-827, -1048) /w:[ 37 -1 38 80 ]
  //: joint g241 (w58) @(195, -1018) /w:[ -1 12 94 11 ]
  _GGOR4 #(10) g5 (.I0(w242), .I1(w240), .I2(w81), .I3(w20), .Z(w88));   //: @(-1068,-562) /sn:0 /R:1 /w:[ 39 33 0 0 1 ]
  _GGAND2 #(6) g118 (.I0(w229), .I1(w155), .Z(w142));   //: @(-506,-939) /sn:0 /w:[ 7 1 1 ]
  _GGCLOCK_P100_0_50 g84 (.Z(w192));   //: @(-1626,-67) /sn:0 /w:[ 103 ] /omega:100 /phi:0 /duty:50
  //: joint g201 (w192) @(-1354, -768) /w:[ 79 80 90 -1 ]
  //: joint g112 (w154) @(-854, -1007) /w:[ 6 -1 5 40 ]
  //: joint g279 (w58) @(195, -827) /w:[ -1 8 98 7 ]
  _GGOR1 #(1) g255 (.I0(w47), .Z(w257));   //: @(82,-1465) /sn:0 /R:1 /w:[ 1 0 ]
  set_flags g21 (.x0_input_01(w95), .x0_input_by_bits(w94), .x0_set_01(w93), .x0_set_by_bits(w24), .x1_input_01(w6), .x1_set_01(w10), .x2_input_01(w35), .x2_input_overflow(w129), .x2_input_parity(w32), .x2_set_01(w35), .x2_set_overflow(w28), .x2_set_parity(w30), .x4_input_01(w36), .x4_input_by_bits(w34), .x4_set_01(w9), .x4_set_by_bits(w207), .x6_input_01(w35), .x6_input_by_bits(w32), .x6_set_01(w35), .x6_set_by_bits(w185), .x7_input_01(w35), .x7_input_by_bits(w32), .x7_set_01(w35), .x7_set_by_bits(w39), .x0_carry_flag(w100), .x0_carry_flag_set(w99), .x1_subtract_flag(w18), .x1_subtract_flag_set(w16), .x2_parity_overflow_flag(w15), .x2_parity_overflow_flag_set(w12), .x4_halfcarry_flag(w8), .x4_halfcarry_flag_set(w2), .x6_zero_flag(w91), .x6_zero_flag_set(w90), .x7_sign_flag(w85), .x7_sign_flag_set(w74));   //: @(629, -904) /sz:(393, 400) /sn:0 /p:[ Li0>1 Li1>3 Li2>3 Li3>0 Li4>0 Li5>0 Li6>19 Li7>0 Li8>11 Li9>15 Li10>3 Li11>3 Li12>1 Li13>1 Li14>3 Li15>3 Li16>11 Li17>9 Li18>7 Li19>3 Li20>3 Li21>5 Li22>0 Li23>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 Ro8<0 Ro9<0 Ro10<0 Ro11<0 ]
  _GGMUX2 #(8, 8) g61 (.I0(w110), .I1(w102), .S(w122), .Z(w116));   //: @(1525,-76) /sn:0 /R:1 /w:[ 0 0 1 0 ] /ss:0 /do:0
  _GGOR9 #(20) g295 (.I0(w93), .I1(w24), .I2(w10), .I3(w28), .I4(w30), .I5(w9), .I6(w207), .I7(w185), .I8(w39), .Z(w111));   //: @(427,-390) /sn:0 /R:3 /w:[ 5 5 5 0 5 0 5 0 0 1 ]
  _GGJKFF #(10, 10, 20) x4_set_b (.Q(w207), ._Q(w208), .J(w209), .K(w237), .PRE(w237), .CLR(w58), .CK(w192));   //: @(158,-611) /w:[ 0 0 1 3 5 103 35 ] /mi:0
  //: joint g32 (w58) @(-961, -1048) /w:[ 39 -1 40 78 ]
  _GGREG8 #(10, 10, 20) g20 (.Q(w144), .D(w145), .EN(w119), .CLR(w58), .CK(w192));   //: @(-1558,-173) /sn:0 /R:1 /w:[ 0 0 1 71 101 ]
  //: joint g311 (w192) @(212, -960) /w:[ -1 17 18 20 ]
  _GGJKFF #(10, 10, 20) x7_set_b (.Q(w39), ._Q(w194), .J(w195), .K(w241), .PRE(w241), .CLR(w58), .CK(w192));   //: @(158,-422) /w:[ 5 0 1 3 5 0 43 ] /mi:0
  //: joint g134 (w242) @(-529, -399) /w:[ 29 30 32 -1 ]
  //: joint g176 (w19) @(-435, -851) /w:[ -1 4 6 3 ]
  assign w25 = w144[2:0]; //: TAP g175 @(-1678,377) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  //: VDD g97 (w239) @(164,-554) /sn:0 /w:[ 0 ]
  //: joint g240 (w58) @(195, -1114) /w:[ -1 14 92 13 ]
  //: joint g148 (w154) @(-714, -1007) /w:[ 12 -1 11 34 ]
  //: joint g15 (w17) @(1527, 121) /w:[ 6 8 5 -1 ]
  //: joint g89 (w32) @(493, -552) /w:[ 4 6 -1 3 ]
  //: joint g252 (w229) @(64, -1093) /w:[ 26 25 -1 28 ]
  //: VDD g247 (w247) @(165,-1317) /sn:0 /w:[ 0 ]
  _GGMUX2x16 #(8, 8) g165 (.I0(w13), .I1(w45), .S(w64), .Z(w14));   //: @(-1678,-1345) /sn:0 /w:[ 0 1 5 0 ] /ss:1 /do:0
  //: joint g147 (w154) @(-587, -1007) /w:[ 16 -1 15 30 ]
  _GGAND2 #(6) g218 (.I0(w139), .I1(w133), .Z(w138));   //: @(-1037,-1279) /sn:0 /R:2 /w:[ 3 7 3 ]
  _GGMUX2x8 #(8, 8) g62 (.I0(w50), .I1(w112), .S(w123), .Z(w87));   //: @(1632,124) /sn:0 /R:2 /w:[ 3 1 1 3 ] /ss:1 /do:0
  //: joint g160 (w192) @(-966, -768) /w:[ 67 68 70 -1 ]
  _GGAND2 #(6) g55 (.I0(w229), .I1(w215), .Z(w53));   //: @(113,-1184) /sn:0 /w:[ 23 1 0 ]
  //: joint g195 (w22) @(-1529, -1521) /w:[ 2 -1 4 1 ]
  _GGJKFF #(10, 10, 20) x2_set_ov (.Q(w28), ._Q(w118), .J(w167), .K(w225), .PRE(w225), .CLR(w58), .CK(w192));   //: @(158,-992) /w:[ 5 0 1 3 5 95 19 ] /mi:0
  //: frame g53 @(557,-1003) /sn:0 /wi:67 /ht:85 /tx:"Unused"
  //: joint g135 (w22) @(-1707, -110) /w:[ -1 6 5 12 ]
  //: joint g139 (w154) @(-1128, -1007) /w:[ 47 -1 48 54 ]
  //: GROUND g13 (w17) @(1446,142) /sn:0 /w:[ 0 ]
  //: joint g308 (w192) @(212, -1346) /w:[ -1 4 6 3 ]
  _GGAND2 #(6) g246 (.I0(w229), .I1(w246), .Z(w197));   //: @(118,-1279) /sn:0 /w:[ 19 1 0 ]
  _GGAND2 #(6) g116 (.I0(w229), .I1(w136), .Z(w135));   //: @(-633,-830) /sn:0 /w:[ 55 1 0 ]
  //: joint g4 (w60) @(-798, -830) /w:[ -1 6 8 5 ]
  //: frame g157 @(-1508,-546) /sn:0 /wi:103 /ht:58 /tx:""
  //: frame g197 @(1436,-115) /sn:0 /wi:235 /ht:365 /tx:"ADD"
  //: joint g271 (w243) @(152, -729) /w:[ -1 1 2 4 ]
  //: joint g17 (w192) @(-1558, -123) /w:[ -1 100 99 102 ]
  //: joint g137 (w27) @(-1095, -1109) /w:[ 5 -1 6 8 ]
  //: joint g280 (w58) @(195, -735) /w:[ -1 6 100 5 ]
  //: joint g282 (w240) @(34, -415) /w:[ -1 17 18 36 ]
  _GGOR1 #(1) g77 (.I0(w240), .Z(w221));   //: @(80,-973) /sn:0 /R:1 /w:[ 7 0 ]
  //: joint g214 (w130) @(-1551, -1342) /w:[ 2 1 8 -1 ]
  //: joint g291 (w240) @(34, -1031) /w:[ 1 2 -1 4 ]
  //: VDD g275 (w232) @(163,-843) /sn:0 /w:[ 0 ]
  //: joint g51 (w35) @(588, -568) /w:[ 2 4 -1 1 ]
  //: GROUND g144 (w46) @(-1613,-1293) /sn:0 /R:1 /w:[ 0 ]
  //: joint g259 (w225) @(153, -1013) /w:[ -1 1 2 4 ]
  //: joint g161 (w192) @(-832, -768) /w:[ 63 64 66 -1 ]
  _GGJKFF #(10, 10, 20) identify_OP (.Q(w59), ._Q(w55), .J(w56), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-1098,-825) /w:[ 9 1 5 55 57 77 73 ] /mi:0
  assign w82 = w13[15:8]; //: TAP g190 @(-1447,-1493) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g296 (w28) @(432, -728) /w:[ 2 -1 4 1 ]
  _GGOR2 #(6) g103 (.I0(w150), .I1(w89), .Z(w163));   //: @(-1439,-1068) /sn:0 /R:2 /w:[ 5 1 0 ]
  _GGOR2 #(6) g65 (.I0(w240), .I1(w242), .Z(w189));   //: @(-412,-728) /sn:0 /R:1 /w:[ 21 0 0 ]
  //: joint g304 (w192) @(212, -489) /w:[ -1 37 38 40 ]
  _GGAND2x8 #(6) g185 (.I0(w50), .I1(w33), .Z(w84));   //: @(294,-251) /sn:0 /R:2 /w:[ 15 5 0 ]
  _GGAND2 #(6) g72 (.I0(w229), .I1(w230), .Z(w187));   //: @(119,-522) /sn:0 /w:[ 51 0 0 ]
  _GGOR1 #(1) g251 (.I0(w242), .Z(w250));   //: @(89,-1359) /sn:0 /R:1 /w:[ 25 0 ]
  _GGJKFF #(10, 10, 20) ADD_DB_DB (.Q(w121), ._Q(w134), .J(w135), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-582,-825) /w:[ 7 0 1 33 31 85 57 ] /mi:0
  _GGOR2 #(6) g6 (.I0(w17), .I1(w17), .Z(w123));   //: @(1560,124) /sn:0 /w:[ 7 3 0 ]
  //: joint g136 (w37) @(-1080, -1104) /w:[ 3 -1 4 6 ]
  //: joint g142 (w1) @(-1311, -1074) /w:[ 2 -1 1 4 ]
  _GGOR1 #(1) g277 (.I0(w242), .Z(w226));   //: @(76,-788) /sn:0 /R:1 /w:[ 15 1 ]
  _GGOR2 #(6) g7 (.I0(w17), .I1(w17), .Z(w122));   //: @(1525,-25) /sn:0 /R:1 /w:[ 13 11 0 ]
  make_negative g58 (.Input0(w50), .Output0(w112));   //: @(1511, 177) /sz:(101, 47) /R:2 /sn:0 /p:[ Bi0>0 To0<0 ]
  //: GROUND g56 (w110) @(1462,-66) /sn:0 /R:3 /w:[ 1 ]
  //: joint g124 (w240) @(-913, -415) /w:[ 27 28 30 -1 ]
  //: joint g297 (w30) @(427, -712) /w:[ 2 -1 1 4 ]
  //: joint g200 (w192) @(-1255, -1243) /w:[ 82 88 81 -1 ]
  //: frame g229 @(1625,-327) /sn:0 /wi:68 /ht:59 /tx:"Overflow"
  //: VDD g98 (w241) @(164,-465) /sn:0 /w:[ 0 ]
  //: joint g204 (w58) @(-1093, -1303) /w:[ 52 -1 51 54 ]
  _GGREG16 #(10, 10, 20) ADDRESS_BUS (.Q(w13), .D(w14), .EN(w46), .CLR(w58), .CK(w192));   //: @(-1678,-1298) /w:[ 11 1 1 59 97 ]
  //: joint g208 (w131) @(-1260, -1315) /w:[ 2 4 -1 1 ]
  //: joint g52 (w35) @(588, -792) /w:[ 18 20 -1 17 ]
  //: joint g40 (w58) @(-1372, -509) /w:[ -1 65 66 68 ]
  _GGOR2 #(6) g81 (.I0(w242), .I1(w240), .Z(w233));   //: @(92,-402) /sn:0 /R:1 /w:[ 27 37 0 ]
  //: joint g313 (w192) @(212, -772) /w:[ -1 25 26 28 ]
  //: joint g108 (w58) @(-451, -1048) /w:[ 31 -1 32 86 ]
  //: joint g210 (w146) @(-964, -1313) /w:[ 2 4 -1 1 ]
  _GGJKFF #(10, 10, 20) x4_set_01 (.Q(w9), ._Q(w214), .J(w210), .K(w243), .PRE(w243), .CLR(w58), .CK(w192));   //: @(157,-707) /w:[ 5 0 1 3 5 101 31 ] /mi:0
  //: joint g131 (w20) @(-1060, -447) /w:[ 2 1 8 -1 ]
  //: joint g299 (w207) @(417, -648) /w:[ 2 -1 1 4 ]
  //: joint g290 (w240) @(34, -949) /w:[ 6 5 -1 8 ]
  //: joint g266 (w58) @(195, -1230) /w:[ -1 16 26 15 ]
  //: SWITCH CLR (CLR) @(-1469,-509) /w:[ 0 ] /st:0 /dn:1
  //: joint g209 (w132) @(-1103, -1317) /w:[ 2 4 -1 1 ]
  //: VDD g96 (w237) @(164,-653) /sn:0 /w:[ 0 ]
  //: joint g294 (w10) @(437, -808) /w:[ 1 -1 2 4 ]
  _GGAND2 #(6) g117 (.I0(w229), .I1(w180), .Z(w128));   //: @(-745,-924) /sn:0 /w:[ 57 1 0 ]
  //: joint g221 (w133) @(-990, -1279) /w:[ 4 3 6 -1 ]
  //: GROUND g315 (w47) @(113,-1434) /sn:0 /R:1 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) DATA_BUS (.Q(w50), .D(w32), .EN(w115), .CLR(~w92), .CK(w192));   //: @(182,-137) /w:[ 19 0 1 1 107 ]
  _GGOR1 #(1) g78 (.I0(w242), .Z(w224));   //: @(77,-882) /sn:0 /R:1 /w:[ 19 1 ]
  _GGOR2 #(6) g155 (.I0(w19), .I1(w121), .Z(w72));   //: @(-473,-832) /sn:0 /w:[ 7 5 0 ]
  //: joint g113 (w154) @(-1103, -1007) /w:[ 45 -1 46 56 ]
  _GGAND2 #(6) g219 (.I0(w139), .I1(w59), .Z(w157));   //: @(-901,-1279) /sn:0 /R:2 /w:[ 0 3 3 ]
  //: joint g223 (w138) @(-1062, -1279) /w:[ 2 -1 4 1 ]
  //: joint g105 (w58) @(-297, -1048) /w:[ 29 -1 30 88 ]
  _GGMUX2x16 #(8, 8) g212 (.I0(w68), .I1(w96), .S(w149), .Z(w45));   //: @(-1609,-1411) /sn:0 /R:3 /w:[ 0 0 1 0 ] /ss:1 /do:0
  //: joint g303 (w192) @(158, -350) /w:[ 41 42 44 -1 ]
  //: joint g292 (w93) @(447, -856) /w:[ 2 -1 1 4 ]
  //: joint g43 (w229) @(-541, -942) /w:[ 6 8 5 -1 ]
  flags g38 (.x0_carry_flag(w100), .x0_change_carry_flag(w99), .x1_change_Subtract_flag(w18), .x1_subtract_flag(w16), .x2_parity_Overflow_flag(w15), .x2_change_Parity_Overflow_flag(w12), .x4_change_Half_carry_flag(w8), .x4_half_carry_flag(w2), .x6_change_zero_flag(w91), .x6_zero_flag(w90), .x7_change_sign_flag(w85), .x7_sign_flag(w74), .Flag_input(w86), .Flag_output(w3));   //: @(1067, -904) /sz:(405, 236) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>1 Li7>1 Li8>1 Li9>1 Li10>1 Li11>1 Bi0>0 Bo0<0 ]
  //: VDD g205 (w131) @(-1249,-1330) /sn:0 /w:[ 5 ]
  //: joint g305 (w192) @(212, -578) /w:[ -1 33 34 36 ]
  //: joint g287 (w242) @(44, -863) /w:[ 18 20 -1 17 ]
  //: joint g48 (w58) @(-704, -1048) /w:[ 35 -1 36 82 ]
  //: joint g276 (w232) @(152, -825) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g237 (.I0(w229), .I1(w235), .Z(w210));   //: @(108,-712) /sn:0 /w:[ 43 1 0 ]
  _GGOR2 #(6) g122 (.I0(w65), .I1(w60), .Z(w229));   //: @(-800,-868) /sn:0 /R:1 /w:[ 0 7 0 ]
  //: joint g95 (w22) @(-1707, -183) /w:[ 8 -1 10 7 ]
  _GGJKFF #(10, 10, 20) addr_2_half (.Q(w130), ._Q(w137), .J(w138), .K(w132), .PRE(w132), .CLR(w58), .CK(w192));   //: @(-1098,-1274) /w:[ 5 0 5 3 0 55 87 ] /mi:1
  _GGOR2 #(6) g80 (.I0(w240), .I1(w242), .Z(w230));   //: @(88,-498) /sn:0 /R:1 /w:[ 15 7 1 ]
  //: joint g170 (w65) @(-938, -924) /w:[ 1 -1 2 4 ]
  _GGMUX2x8 #(8, 8) g178 (.I0(w11), .I1(w41), .S(w76), .Z(w32));   //: @(182,-229) /sn:0 /w:[ 0 1 1 13 ] /ss:0 /do:0
  assign w23 = w13[7:0]; //: TAP g189 @(-1538,-1493) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g182 (w121) @(-149, -298) /w:[ 1 2 -1 8 ]
  //: joint g269 (w229) @(64, -619) /w:[ 46 45 -1 48 ]
  //: VDD g90 (w26) @(164,-1218) /sn:0 /w:[ 0 ]
  _GGOR4 #(10) g128 (.I0(w37), .I1(w27), .I2(w157), .I3(w138), .Z(w89));   //: @(-1145,-1111) /sn:0 /R:2 /w:[ 5 7 0 0 0 ]
  assign w143 = w144[5:3]; //: TAP g174 @(-1678,294) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  instruction_decoder g2 (.Instruction_input(w144), .LD_r_r(w20), .LD_r_n(w81), .ADD_A_n(w240), .AND_A_n(w242), .JP_nn(w38), .NOP(w48));   //: @(-1399, -463) /sz:(247, 587) /sn:0 /p:[ Li0>3 Ro0<9 Ro1<9 Ro2<35 Ro3<41 Ro4<1 Ro5<0 ]
  //: joint g268 (w58) @(195, -1405) /w:[ -1 20 22 19 ]
  //: joint g91 (w192) @(-1594, -768) /w:[ 91 92 -1 98 ]
  //: joint g141 (w58) @(-1207, -1048) /w:[ 43 -1 44 74 ]
  //: joint g265 (w229) @(64, -906) /w:[ 34 33 -1 36 ]
  //: joint g285 (w242) @(44, -654) /w:[ 10 12 -1 9 ]
  //: joint g29 (w154) @(-327, -1007) /w:[ 22 -1 21 24 ]
  //: joint g288 (w242) @(44, -1045) /w:[ 22 24 -1 21 ]
  //: joint g168 (w50) @(182, -35) /w:[ 10 12 -1 9 ]
  //: joint g278 (w229) @(64, -812) /w:[ 38 37 -1 40 ]
  _GGOR1 #(1) g18 (.I0(w20), .Z(w70));   //: @(-1024,-875) /sn:0 /R:1 /w:[ 7 0 ]
  //: joint g199 (w192) @(-1098, -1243) /w:[ 84 86 83 -1 ]
  _GGAND2 #(6) g119 (.I0(w72), .I1(w189), .Z(w152));   //: @(-395,-830) /sn:0 /w:[ 1 1 0 ]
  //: joint g173 (w144) @(-1676, -112) /w:[ 5 6 -1 8 ]
  //: joint g154 (w229) @(-788, -896) /w:[ 4 -1 3 54 ]
  //: joint g256 (w229) @(64, -1000) /w:[ 30 29 -1 32 ]
  //: joint g188 (w13) @(-1736, -1376) /w:[ 1 2 -1 8 ]
  //: joint g184 (w50) @(182, -93) /w:[ 14 16 -1 13 ]
  //: joint g172 (w60) @(-161, -189) /w:[ 1 2 -1 12 ]
  //: joint g50 (w229) @(64, -1282) /w:[ 18 17 -1 20 ]
  //: joint g261 (w231) @(153, -919) /w:[ -1 1 2 4 ]
  //: joint g193 (w50) @(1642, 234) /w:[ -1 2 1 4 ]
  _GGAND2 #(6) g73 (.I0(w229), .I1(w233), .Z(w195));   //: @(117,-427) /sn:0 /w:[ 53 1 0 ]
  //: SWITCH g9 (w92) @(244,-182) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g102 (w35) @(588, -600) /w:[ 6 8 -1 5 ]
  //: joint g186 (w33) @(963, 46) /w:[ 3 4 6 -1 ]
  _GGAND2 #(6) g71 (.I0(w229), .I1(w227), .Z(w209));   //: @(109,-616) /sn:0 /w:[ 47 1 0 ]
  _GGADD8 #(68, 70, 62, 64) g59 (.A(w87), .B(w33), .S(w29), .CI(w116), .CO(w94));   //: @(1616,0) /sn:0 /R:2 /w:[ 0 0 0 5 5 ]
  _GGAND2 #(6) g169 (.I0(w60), .I1(!w65), .Z(w124));   //: @(-9,-100) /sn:0 /w:[ 13 9 0 ]
  //: joint g249 (w229) @(64, -1187) /w:[ 22 21 -1 24 ]
  //: GROUND g99 (w35) @(588,-974) /sn:0 /R:2 /w:[ 21 ]
  _GGMUX2x8 #(8, 8) g180 (.I0(w29), .I1(w84), .S(w125), .Z(w41));   //: @(247,-261) /sn:0 /R:3 /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: joint g45 (w31) @(-1861, -1102) /w:[ 2 1 -1 4 ]
  //: joint g36 (w154) @(-1197, -1007) /w:[ 49 50 -1 52 ]
  _GGJKFF #(10, 10, 20) x1_set_01 (.Q(w10), ._Q(w78), .J(w79), .K(w219), .PRE(w219), .CLR(w58), .CK(w192));   //: @(158,-1085) /w:[ 3 0 1 3 5 93 15 ] /mi:0
  _GGADD16 #(132, 134, 126, 128) g69 (.A(w31), .B(w168), .S(w158), .CI(w166), .CO(w182));   //: @(-1528,-1132) /sn:0 /w:[ 0 1 0 1 0 ]
  //: joint g156 (w58) @(-1372, -1048) /w:[ 45 46 -1 60 ]
  _GGAND2 #(6) g254 (.I0(w229), .I1(w257), .Z(w5));   //: @(107,-1490) /sn:0 /w:[ 11 1 0 ]
  //: joint g273 (w240) @(-414, -415) /w:[ 19 20 22 -1 ]
  //: joint g191 (w86) @(1322, -546) /w:[ 2 1 -1 4 ]
  assign w67 = w33[3:0]; //: TAP g232 @(1570,44) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w61 = w87[3:0]; //: TAP g233 @(1630,81) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  _GGOR1 #(1) g239 (.I0(w242), .Z(w235));   //: @(82,-682) /sn:0 /R:1 /w:[ 11 0 ]
  _GGOR1 #(1) g28 (.I0(w242), .Z(w155));   //: @(-529,-814) /sn:0 /R:1 /w:[ 31 0 ]
  _GGAND2 #(6) g57 (.I0(w229), .I1(w218), .Z(w79));   //: @(111,-1090) /sn:0 /w:[ 27 1 0 ]
  //: joint g242 (w58) @(195, -921) /w:[ -1 10 96 9 ]
  _GGJKFF #(10, 10, 20) x0_set_01 (.Q(w93), ._Q(w252), .J(w211), .K(w254), .PRE(w254), .CLR(w58), .CK(w192));   //: @(155,-1379) /w:[ 0 0 1 3 5 23 7 ] /mi:0
  //: joint g286 (w242) @(44, -762) /w:[ 14 16 -1 13 ]
  _GGNOR3 #(6) g150 (.I0(w60), .I1(w56), .I2(w64), .Z(w4));   //: @(-1718,-666) /sn:0 /R:2 /w:[ 11 0 0 0 ]
  _GGMUX2x8 #(8, 8) g11 (.I0(w144), .I1(w22), .S(w56), .Z(w145));   //: @(-1635,-173) /sn:0 /R:1 /w:[ 7 9 9 1 ] /ss:1 /do:0
  //: joint g14 (w17) @(1511, 126) /w:[ 2 4 1 -1 ]
  //: joint g123 (w229) @(-800, -896) /w:[ 2 56 -1 1 ]
  //: joint g187 (w192) @(-188, -137) /w:[ 106 105 -1 108 ]
  _GGROM16x8 #(10, 30) instructions_rom (.A(w31), .D(w22), .OE(w4));   //: @(-1752,-182) /w:[ 9 11 1 ] /mem:"/home/pawel/Desktop/OIAK/oiak-projekt/instructions.mem"
  _GGOR1 #(1) g79 (.I0(w240), .Z(w227));   //: @(83,-586) /sn:0 /R:1 /w:[ 11 0 ]
  _GGAND2 #(6) g115 (.I0(w59), .I1(w175), .Z(w150));   //: @(-901,-830) /sn:0 /w:[ 7 1 0 ]
  //: joint g145 (w192) @(-1594, -887) /w:[ 94 -1 96 93 ]
  //: frame g235 @(1682,-62) /sn:0 /wi:132 /ht:108 /tx:"Half_Carry"
  //: joint g236 (w35) @(588, -632) /w:[ 10 12 -1 9 ]
  //: joint g129 (w37) @(-685, -924) /w:[ -1 2 8 1 ]
  _GGOR1 #(1) g27 (.I0(w240), .Z(w136));   //: @(-660,-711) /sn:0 /R:1 /w:[ 25 0 ]
  //: joint g202 (w58) @(-1372, -1303) /w:[ 48 -1 58 47 ]
  //: joint g227 (w63) @(-1297, -1279) /w:[ 2 -1 4 1 ]
  //: joint g171 (w65) @(-175, -184) /w:[ 6 5 -1 8 ]
  _GGJKFF #(10, 10, 20) n_DB (.Q(w60), ._Q(w113), .J(w150), .K(w154), .PRE(w154), .CLR(w58), .CK(w192));   //: @(-832,-825) /w:[ 9 0 3 41 39 81 65 ] /mi:0
  //: VDD g238 (w243) @(163,-749) /sn:0 /w:[ 0 ]
  //: joint g88 (w32) @(182, -159) /w:[ 2 12 -1 1 ]
  //: GROUND g314 (w43) @(112,-1132) /sn:0 /R:1 /w:[ 0 ]
  //: joint g140 (w58) @(-1093, -1048) /w:[ 41 -1 42 76 ]
  //: VDD g207 (w146) @(-953,-1330) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin instruction_decoder
module instruction_decoder(AND_A_n, NOP, JP_nn, ADD_A_n, LD_r_n, LD_r_r, Instruction_input);
//: interface  /sz:(247, 587) /bd:[ Li0>Instruction_input[7:0](16/587) Ro0<LD_r_r(16/587) Ro1<LD_r_n(32/587) Ro2<ADD_A_n(48/587) Ro3<AND_A_n(64/587) Ro4<JP_nn(80/587) Ro5<NOP(96/587) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output ADD_A_n;    //: /sn:0 {0}(654,687)(654,306){1}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
output NOP;    //: /sn:0 {0}(1847,587)(1847,324)(1752,324)(1752,306){1}
output AND_A_n;    //: /sn:0 {0}(464,633)(464,306){1}
supply1 w127;    //: /sn:0 {0}(1090,400)(1090,437){1}
//: {2}(1092,439)(1132,439){3}
//: {4}(1136,439)(1152,439){5}
//: {6}(1156,439)(1172,439){7}
//: {8}(1176,439)(1194,439)(1194,469){9}
//: {10}(1174,441)(1174,469){11}
//: {12}(1154,441)(1154,469){13}
//: {14}(1134,441)(1134,469){15}
//: {16}(1090,441)(1090,456)(1114,456)(1114,469){17}
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
output LD_r_n;    //: /sn:0 {0}(1624,513)(1624,473){1}
output LD_r_r;    //: /sn:0 {0}(1313,481)(1313,444){1}
output JP_nn;    //: /sn:0 {0}(706,535)(706,466)(664,466)(664,306){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire HALT;    //: /sn:0 {0}(1156,562)(1156,580)(1276,580)(1276,365)(1292,365)(1292,378){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire ED;    //: /sn:0 {0}(-39,539)(439,539)(439,306){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w109;    //: /sn:0 {0}(989,160)(989,394){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w19;    //: /sn:0 {0}(633,317)(633,306){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w54;    //: /sn:0 {0}(1139,469)(1139,339)(1227,339)(1227,317){1}
wire w91;    //: /sn:0 {0}(1161,541)(1161,505)(1176,505)(1176,490){1}
wire w86;    //: /sn:0 {0}(1179,469)(1179,379)(1247,379)(1247,317){1}
wire CPL_negation;    //: /sn:0 {0}(1539,306)(1539,615){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire DD;    //: /sn:0 {0}(-52,560)(540,560)(540,306){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,397)(1609,397)(1609,452){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w8;    //: /sn:0 {0}(1310,423)(1310,207)(254,207){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w260;    //: /sn:0 {0}(1619,452)(1619,375)(1571,375)(1571,306){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire ADD_A_r;    //: /sn:0 {0}(1006,458)(1006,435)(1006,435)(1006,415){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w11;    //: /sn:0 {0}(944,394)(944,314){1}
//: {2}(946,312)(964,312)(964,394){3}
//: {4}(944,310)(944,218)(254,218){5}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,391)(1639,391)(1639,452){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w55;    //: /sn:0 {0}(969,160)(969,394){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire SBC_A_r;    //: /sn:0 {0}(939,511)(939,461)(946,461)(946,415){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w286;    //: /sn:0 {0}(1624,452)(1624,306){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w6;    //: /sn:0 {0}(1320,423)(1320,200)(254,200){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w7;    //: /sn:0 {0}(1315,423)(1315,204)(254,204){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire FD;    //: /sn:0 {0}(-41,487)(343,487)(343,306){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w72;    //: /sn:0 {0}(1237,317)(1237,364)(1159,364)(1159,469){1}
wire w278;    //: /sn:0 {0}(1629,452)(1629,375)(1652,375)(1652,306){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w36;    //: /sn:0 {0}(1305,423)(1305,414)(1294,414)(1294,399){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w10;    //: /sn:0 {0}(1004,394)(1004,312)(986,312){1}
//: {2}(984,310)(984,214)(254,214){3}
//: {4}(984,314)(984,394){5}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire SUB_r;    //: /sn:0 {0}(966,458)(966,437)(966,437)(966,415){1}
wire CB;    //: /sn:0 {0}(636,306)(636,582)(-15,582){1}
wire w130;    //: /sn:0 {0}(1009,160)(1009,394){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w108;    //: /sn:0 {0}(1199,469)(1199,412)(1257,412)(1257,317){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(948,156){13}
//: {14}(949,156)(968,156){15}
//: {16}(969,156)(988,156){17}
//: {18}(989,156)(1008,156){19}
//: {20}(1009,156)(1240,156){21}
//: {22}(1244,156)(1481,156){23}
//: {24}(#:1485,156)(1564,156){25}
//: {26}(#:1568,156)(1645,156){27}
//: {28}(#:1649,156)(1726,156)(1726,277){29}
//: {30}(1647,158)(1647,277){31}
//: {32}(1566,158)(1566,277){33}
//: {34}(1483,158)(1483,277){35}
//: {36}(1242,158)(#:1242,311){37}
//: {38}(842,158)(842,277){39}
//: {40}(744,158)(744,277){41}
//: {42}(649,158)(649,277){43}
//: {44}(560,158)(560,277){45}
//: {46}(459,158)(459,277){47}
//: {48}(363,158)(363,277){49}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w268;    //: /sn:0 {0}(1614,452)(1614,389)(1543,389)(1543,306){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w304;    //: /sn:0 {0}(1634,452)(1634,381)(1703,381)(1703,306){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w33;    //: /sn:0 {0}(949,160)(949,394){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w69;    //: /sn:0 {0}(1151,541)(1151,505)(1136,505)(1136,490){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w277;    //: /sn:0 {0}(1655,328)(1655,306){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire OR_A_n;    //: /sn:0 {0}(368,637)(368,306){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w85;    //: /sn:0 {0}(1156,541)(1156,490){1}
wire w126;    //: /sn:0 {0}(1196,490)(1196,526)(1166,526)(1166,541){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire ADC_A_r;    //: /sn:0 {0}(986,511)(986,462)(986,462)(986,415){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w9;    //: /sn:0 {0}(1297,378)(1297,290)(1086,290){1}
//: {2}(1084,288)(1084,211)(254,211){3}
//: {4}(1084,292)(1084,380)(1119,380)(1119,469){5}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w51;    //: /sn:0 {0}(1116,490)(1116,526)(1146,526)(1146,541){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire XOR_A_n;    //: /sn:0 {0}(436,660)(436,306){1}
//: enddecls

  //: joint g44 (w127) @(1134, 439) /w:[ 4 -1 3 14 ]
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(OR_A_n), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(FD), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g47 (w9) @(1084, 290) /w:[ 1 2 -1 4 ]
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(CPL_negation));   //: @(1566,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 ] /ss:0 /do:1
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 38 ]
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  _GGAND2 #(6) g30 (.I0(w108), .I1(!w127), .Z(w126));   //: @(1196,480) /sn:0 /R:3 /w:[ 0 9 0 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 44 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 1 1 1 3 3 5 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 42 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  assign w130 = w1[3]; //: TAP g60 @(1009,154) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  _GGAND2 #(6) g29 (.I0(w86), .I1(w127), .Z(w91));   //: @(1176,480) /sn:0 /R:3 /w:[ 0 11 1 ]
  //: OUT g70 (AND_A_n) @(464,630) /sn:0 /R:3 /w:[ 0 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 31 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 ] /ss:0 /do:1
  _GGAND2 #(6) g10 (.I0(w33), .I1(w11), .Z(SBC_A_r));   //: @(946,405) /sn:0 /R:3 /w:[ 1 0 1 ]
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 40 ]
  _GGAND2 #(6) g65 (.I0(w9), .I1(!HALT), .Z(w36));   //: @(1294,389) /sn:0 /R:3 /w:[ 0 1 1 ]
  assign {w54, w72, w86, w108} = w1; //: CONCAT g49  @(1242,312) /sn:0 /R:1 /w:[ 1 0 1 1 37 ] /dr:0 /tp:0 /drp:0
  _GGAND5 #(12) g50 (.I0(w126), .I1(w91), .I2(w85), .I3(w69), .I4(w51), .Z(HALT));   //: @(1156,552) /sn:0 /R:3 /w:[ 1 0 0 0 1 0 ]
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(DD), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 ] /ss:0 /do:1
  //: OUT g68 (NOP) @(1847,584) /sn:0 /R:3 /w:[ 0 ]
  assign w55 = w1[3]; //: TAP g58 @(969,154) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: joint g56 (w10) @(984, 312) /w:[ 1 2 -1 4 ]
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(JP_nn), .Z4(w78), .Z5(w79), .Z6(ADD_A_n), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(CB), .Z12(w19), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 43 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 28 -1 27 30 ]
  //: OUT g73 (JP_nn) @(706,532) /sn:0 /R:3 /w:[ 0 ]
  assign w109 = w1[3]; //: TAP g59 @(989,154) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  //: VDD g31 (w127) @(1101,400) /sn:0 /w:[ 0 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 46 ]
  //: OUT g67 (ADD_A_n) @(654,684) /sn:0 /R:3 /w:[ 0 ]
  //: joint g45 (w127) @(1154, 439) /w:[ 6 -1 5 12 ]
  //: joint g33 (w1) @(1483, 156) /w:[ 24 -1 23 34 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: OUT g54 (LD_r_n) @(1624,510) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g52 (LD_r_r) @(1313,478) /sn:0 /R:3 /w:[ 0 ]
  _GGOR4 #(10) g12 (.I0(w6), .I1(w7), .I2(w8), .I3(w36), .Z(LD_r_r));   //: @(1313,434) /sn:0 /R:3 /w:[ 0 0 0 0 1 ]
  assign w33 = w1[3]; //: TAP g57 @(949,154) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  _GGAND2 #(6) g28 (.I0(!w130), .I1(w10), .Z(ADD_A_r));   //: @(1006,405) /sn:0 /R:3 /w:[ 1 0 1 ]
  //: joint g46 (w127) @(1174, 439) /w:[ 8 -1 7 10 ]
  //: joint g34 (w1) @(1566, 156) /w:[ 26 -1 25 32 ]
  _GGAND2 #(6) g11 (.I0(!w55), .I1(w11), .Z(SUB_r));   //: @(966,405) /sn:0 /R:3 /w:[ 1 3 1 ]
  _GGAND2 #(6) g14 (.I0(w54), .I1(!w127), .Z(w69));   //: @(1136,480) /sn:0 /R:3 /w:[ 0 15 1 ]
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(AND_A_n), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(ED), .Z14(XOR_A_n), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(NOP), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 29 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 48 ]
  //: joint g32 (w127) @(1090, 439) /w:[ 2 1 -1 16 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  _GGAND2 #(6) g15 (.I0(w72), .I1(w127), .Z(w85));   //: @(1156,480) /sn:0 /R:3 /w:[ 1 13 1 ]
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGAND2 #(6) g27 (.I0(w109), .I1(w10), .Z(ADC_A_r));   //: @(986,405) /sn:0 /R:3 /w:[ 1 5 1 ]
  //: joint g48 (w1) @(1242, 156) /w:[ 22 -1 21 36 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  //: joint g55 (w11) @(944, 312) /w:[ 2 4 -1 1 ]
  _GGAND2 #(6) g13 (.I0(w9), .I1(w127), .Z(w51));   //: @(1116,480) /sn:0 /R:3 /w:[ 5 17 0 ]
  _GGOR7 #(16) g53 (.I0(w296), .I1(w304), .I2(w278), .I3(w286), .I4(w260), .I5(w268), .I6(w250), .Z(LD_r_n));   //: @(1624,463) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin instruction_IY
module instruction_IY(CB, Instruction_input);
//: interface  /sz:(303, 511) /bd:[ Li0>Instruction_input[7:0](204/511) Bo0<CB(20/303) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
output CB;    //: /sn:0 {0}(-67,486)(636,486)(636,306){1}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire w139;    //: /sn:0 {0}(924,306)(924,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire w128;    //: /sn:0 {0}(963,306)(963,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w86;    //: /sn:0 {0}(633,306)(633,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,321){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w140;    //: /sn:0 {0}(921,306)(921,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w147;    //: /sn:0 {0}(1049,306)(1049,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w260;    //: /sn:0 {0}(1571,306)(1571,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w44;    //: /sn:0 {0}(464,306)(464,321){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w135;    //: /sn:0 {0}(938,306)(938,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w11;    //: /sn:0 {0}(254,218)(898,218)(898,290)(913,290){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,321){1}
wire w129;    //: /sn:0 {0}(959,306)(959,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w286;    //: /sn:0 {0}(1624,306)(1624,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w158;    //: /sn:0 {0}(1011,306)(1011,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w142;    //: /sn:0 {0}(914,306)(914,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w148;    //: /sn:0 {0}(1046,306)(1046,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w154;    //: /sn:0 {0}(1025,306)(1025,321){1}
wire w156;    //: /sn:0 {0}(1018,306)(1018,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w130;    //: /sn:0 {0}(956,306)(956,321){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w131;    //: /sn:0 {0}(952,306)(952,321){1}
wire w268;    //: /sn:0 {0}(1543,306)(1543,321){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w304;    //: /sn:0 {0}(1703,306)(1703,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w52;    //: /sn:0 {0}(436,306)(436,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w150;    //: /sn:0 {0}(1039,306)(1039,321){1}
wire w33;    //: /sn:0 {0}(343,306)(343,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w69;    //: /sn:0 {0}(540,306)(540,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w146;    //: /sn:0 {0}(1053,306)(1053,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w151;    //: /sn:0 {0}(1035,306)(1035,321){1}
wire w161;    //: /sn:0 {0}(1000,306)(1000,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w137;    //: /sn:0 {0}(931,306)(931,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w157;    //: /sn:0 {0}(1014,306)(1014,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w132;    //: /sn:0 {0}(949,306)(949,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w152;    //: /sn:0 {0}(1032,306)(1032,321){1}
wire w138;    //: /sn:0 {0}(928,306)(928,321){1}
wire w269;    //: /sn:0 {0}(1539,306)(1539,321){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w136;    //: /sn:0 {0}(935,306)(935,321){1}
wire w134;    //: /sn:0 {0}(942,306)(942,321){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w153;    //: /sn:0 {0}(1028,306)(1028,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w155;    //: /sn:0 {0}(1021,306)(1021,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w26;    //: /sn:0 {0}(368,306)(368,321){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w143;    //: /sn:0 {0}(910,306)(910,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w278;    //: /sn:0 {0}(1652,306)(1652,321){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w159;    //: /sn:0 {0}(1007,306)(1007,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w141;    //: /sn:0 {0}(917,306)(917,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w10;    //: /sn:0 {0}(254,214)(988,214)(988,290)(1003,290){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(935,156){13}
//: {14}(#:939,156)(1025,156){15}
//: {16}(#:1029,156)(1118,156){17}
//: {18}(#:1122,156)(1208,156){19}
//: {20}(#:1212,156)(1297,156){21}
//: {22}(#:1301,156)(1391,156){23}
//: {24}(#:1395,156)(1481,156){25}
//: {26}(#:1485,156)(1564,156){27}
//: {28}(#:1568,156)(1645,156){29}
//: {30}(#:1649,156)(1726,156)(1726,277){31}
//: {32}(1647,158)(1647,277){33}
//: {34}(1566,158)(1566,277){35}
//: {36}(1483,158)(1483,277){37}
//: {38}(1393,158)(1393,277){39}
//: {40}(1299,158)(1299,277){41}
//: {42}(1210,158)(1210,277){43}
//: {44}(1120,158)(1120,277){45}
//: {46}(1027,158)(1027,277){47}
//: {48}(937,158)(937,277){49}
//: {50}(842,158)(842,277){51}
//: {52}(744,158)(744,277){53}
//: {54}(649,158)(649,277){55}
//: {56}(560,158)(560,277){57}
//: {58}(459,158)(459,277){59}
//: {60}(363,158)(363,277){61}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w290;    //: /sn:0 {0}(1752,306)(1752,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w80;    //: /sn:0 {0}(654,306)(654,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire w277;    //: /sn:0 {0}(1655,306)(1655,321){1}
wire w149;    //: /sn:0 {0}(1042,306)(1042,321){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w160;    //: /sn:0 {0}(1004,306)(1004,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire w133;    //: /sn:0 {0}(945,306)(945,321){1}
wire w77;    //: /sn:0 {0}(664,306)(664,321){1}
wire w51;    //: /sn:0 {0}(439,306)(439,321){1}
//: enddecls

  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 53 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(w26), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(w33), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 61 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 37 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 50 ]
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(w269));   //: @(1566,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w1) @(1210, 156) /w:[ 20 -1 19 42 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 56 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 54 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g29 (w1) @(1120, 156) /w:[ 18 -1 17 44 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 52 ]
  _GGDECODER16 #(6, 6) g10 (.I(w1), .E(w11), .Z0(w128), .Z1(w129), .Z2(w130), .Z3(w131), .Z4(w132), .Z5(w133), .Z6(w134), .Z7(w135), .Z8(w136), .Z9(w137), .Z10(w138), .Z11(w139), .Z12(w140), .Z13(w141), .Z14(w142), .Z15(w143));   //: @(937,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(w69), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 57 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 30 -1 29 32 ]
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 51 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(w77), .Z4(w78), .Z5(w79), .Z6(w80), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(CB), .Z12(w86), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 55 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w1) @(1299, 156) /w:[ 22 -1 21 40 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 58 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: joint g33 (w1) @(1483, 156) /w:[ 26 -1 25 36 ]
  //: OUT g40 (CB) @(-64,486) /sn:0 /R:2 /w:[ 0 ]
  _GGDECODER16 #(6, 6) g12 (.I(w1), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g34 (w1) @(1566, 156) /w:[ 28 -1 27 34 ]
  //: joint g28 (w1) @(1027, 156) /w:[ 16 -1 15 46 ]
  _GGDECODER16 #(6, 6) g14 (.I(w1), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g11 (.I(w1), .E(w10), .Z0(w146), .Z1(w147), .Z2(w148), .Z3(w149), .Z4(w150), .Z5(w151), .Z6(w152), .Z7(w153), .Z8(w154), .Z9(w155), .Z10(w156), .Z11(w157), .Z12(w158), .Z13(w159), .Z14(w160), .Z15(w161));   //: @(1027,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(w44), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(w51), .Z14(w52), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 59 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 60 ]
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(w290), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 31 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g32 (w1) @(1393, 156) /w:[ 24 -1 23 38 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w1), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: joint g27 (w1) @(937, 156) /w:[ 14 -1 13 48 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w1), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 43 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin flags_status
module flags_status(Flag_2_parity_overflow, Flag_1_substract, Flag_0_carry, Flag_6_zero, Flag_7_sign, Flag_4_halfcarry, flags_in);
//: interface  /sz:(351, 112) /bd:[ Li0>flags_in[7:0](16/112) Ro0<Flag_7_sign(96/112) Ro1<Flag_6_zero(80/112) Ro2<Flag_4_halfcarry(64/112) Ro3<Flag_2_parity_overflow(48/112) Ro4<Flag_1_substract(32/112) Ro5<Flag_0_carry(16/112) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Flag_1_substract;    //: /sn:0 {0}(640,148)(396,148){1}
output Flag_6_zero;    //: /sn:0 {0}(640,198)(517,198)(517,198)(396,198){1}
output Flag_0_carry;    //: /sn:0 {0}(640,138)(517,138)(517,138)(396,138){1}
output Flag_2_parity_overflow;    //: /sn:0 {0}(640,158)(519,158)(519,158)(396,158){1}
output Flag_4_halfcarry;    //: /sn:0 {0}(640,178)(518,178)(518,178)(396,178){1}
input [7:0] flags_in;    //: /sn:0 {0}(#:390,173)(#:316,173){1}
output Flag_7_sign;    //: /sn:0 {0}(640,208)(517,208)(517,208)(396,208){1}
wire w3;    //: /sn:0 {0}(396,168)(492,168)(492,99){1}
wire w5;    //: /sn:0 {0}(529,95)(529,188)(396,188){1}
//: enddecls

  //: LED g8 (w3) @(492,92) /sn:0 /w:[ 1 ] /type:0
  //: OUT g4 (Flag_2_parity_overflow) @(637,158) /sn:0 /w:[ 0 ]
  //: OUT g3 (Flag_1_substract) @(637,148) /sn:0 /w:[ 0 ]
  //: OUT g2 (Flag_0_carry) @(637,138) /sn:0 /w:[ 0 ]
  assign {Flag_7_sign, Flag_6_zero, w5, Flag_4_halfcarry, w3, Flag_2_parity_overflow, Flag_1_substract, Flag_0_carry} = flags_in; //: CONCAT g1  @(391,173) /sn:0 /R:2 /w:[ 1 1 1 1 0 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  //: OUT g6 (Flag_6_zero) @(637,198) /sn:0 /w:[ 0 ]
  //: LED g9 (w5) @(529,88) /sn:0 /w:[ 0 ] /type:0
  //: OUT g7 (Flag_7_sign) @(637,208) /sn:0 /w:[ 0 ]
  //: OUT g5 (Flag_4_halfcarry) @(637,178) /sn:0 /w:[ 0 ]
  //: IN g0 (flags_in) @(314,173) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin registers
module registers(Accumulator_input, Flag_input_choose, Clock, _CLR, Register_output1, Register_input_choose, Register_output_choose1, Register_input_dec, Register_input, Accumulator_output, Flag_output, Accumulator_input_choose, Flag_input);
//: interface  /sz:(357, 455) /bd:[ Li0>Accumulator_input[7:0](41/455) Li1>Accumulator_input_choose(82/455) Li2>Clock(124/455) Li3>Flag_input[7:0](165/455) Li4>Flag_input_choose(206/455) Li5>Register_input[7:0](248/455) Li6>Register_input_choose[2:0](289/455) Li7>Register_input_dec(330/455) Li8>Register_output_choose1[2:0](372/455) Li9>_CLR(413/455) Ro0<Accumulator_output[7:0](41/455) Ro1<Flag_output[7:0](82/455) Ro2<Register_output1[7:0](124/455) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Register_input;    //: /sn:0 {0}(#:132,301)(46,301){1}
//: {2}(44,299)(44,267)(382,267){3}
//: {4}(42,301)(-338,301){5}
//: {6}(-340,299)(-340,-50){7}
//: {8}(-338,-52)(244,-52){9}
//: {10}(248,-52)(491,-52)(#:491,-10){11}
//: {12}(246,-50)(246,-17){13}
//: {14}(-342,-52)(-452,-52)(-452,-52)(#:-501,-52){15}
//: {16}(-340,303)(-340,507){17}
//: {18}(-338,509)(-54,509){19}
//: {20}(-50,509)(119,509){21}
//: {22}(-52,507)(-52,474)(382,474){23}
//: {24}(#:-340,511)(-340,707)(21,707){25}
//: {26}(25,707)(122,707){27}
//: {28}(23,705)(23,666)(383,666){29}
supply0 w58;    //: /sn:0 {0}(280,545)(266,545){1}
supply0 w59;    //: /sn:0 {0}(518,545)(511,545){1}
output [7:0] Register_output1;    //: /sn:0 {0}(#:2161,425)(2344,425)(2344,425)(#:2515,425){1}
input [2:0] Register_input_choose;    //: /sn:0 {0}(#:-501,-118)(#:-257,-118){1}
input Accumulator_input_choose;    //: /sn:0 {0}(118,32)(118,3){1}
//: {2}(120,1)(164,1){3}
//: {4}(118,-1)(118,-651){5}
supply0 w60;    //: /sn:0 {0}(289,742)(266,742){1}
input Clock;    //: /sn:0 {0}(190,540)(173,540){1}
//: {2}(171,538)(171,427){3}
//: {4}(173,425)(423,425){5}
//: {6}(425,423)(425,335){7}
//: {8}(427,333)(435,333){9}
//: {10}(425,331)(425,156)(434,156){11}
//: {12}(425,427)(425,538){13}
//: {14}(427,540)(435,540){15}
//: {16}(425,542)(425,737)(435,737){17}
//: {18}(171,423)(171,335){19}
//: {20}(173,333)(190,333){21}
//: {22}(171,331)(171,158){23}
//: {24}(173,156)(189,156){25}
//: {26}(169,156)(60,156)(60,-266)(-97,-266){27}
//: {28}(171,542)(171,737)(190,737){29}
input Register_input_dec;    //: /sn:0 {0}(-501,-216)(-246,-216){1}
//: {2}(-242,-216)(139,-216)(139,-4)(164,-4){3}
//: {4}(-244,-214)(-244,-142){5}
input [7:0] Flag_input;    //: /sn:0 {0}(#:471,-10)(471,-475)(567,-475)(#:567,-488){1}
output [7:0] Accumulator_output;    //: /sn:0 {0}(216,63)(216,47)(#:157,47)(157,217)(224,217){1}
//: {2}(228,217)(318,217){3}
//: {4}(322,217)(#:1627,217)(1627,448)(#:2132,448){5}
//: {6}(320,215)(320,-218)(320,-218)(320,-656){7}
//: {8}(226,215)(#:226,167){9}
supply0 w54;    //: /sn:0 {0}(540,161)(510,161){1}
output [7:0] Flag_output;    //: /sn:0 {0}(#:655,-651)(655,-443)(531,-443)(531,204)(473,204){1}
//: {2}(471,202)(#:471,167){3}
//: {4}(469,204)(410,204)(410,53)(461,53)(461,78){5}
supply0 w52;    //: /sn:0 {0}(281,161)(265,161){1}
input _CLR;    //: /sn:0 {0}(510,151)(558,151){1}
//: {2}(560,149)(560,-300)(339,-300){3}
//: {4}(335,-300)(-64,-300){5}
//: {6}(337,-298)(337,149){7}
//: {8}(335,151)(265,151){9}
//: {10}(337,153)(337,326){11}
//: {12}(335,328)(266,328){13}
//: {14}(337,330)(337,533){15}
//: {16}(335,535)(266,535){17}
//: {18}(337,537)(337,732)(266,732){19}
//: {20}(560,153)(560,326){21}
//: {22}(558,328)(511,328){23}
//: {24}(560,330)(560,533){25}
//: {26}(558,535)(511,535){27}
//: {28}(560,537)(560,732)(511,732){29}
input [2:0] Register_output_choose1;    //: /sn:0 {0}(#:2086,-150)(2148,-150)(2148,402){1}
input [7:0] Accumulator_input;    //: /sn:0 {0}(226,-17)(226,-209)(226,-209)(#:226,-401){1}
supply0 w55;    //: /sn:0 {0}(285,338)(266,338){1}
supply0 w61;    //: /sn:0 {0}(525,742)(511,742){1}
input Flag_input_choose;    //: /sn:0 {0}(480,-651)(480,-497)(421,-497)(421,4){1}
//: {2}(423,6)(458,6){3}
//: {4}(421,8)(421,94)(448,94){5}
supply0 w57;    //: /sn:0 {0}(534,338)(511,338){1}
wire [7:0] w13;    //: /sn:0 {0}(#:472,344)(472,389){1}
//: {2}(474,391)(#:1553,391)(1553,408)(#:2132,408){3}
//: {4}(470,391)(#:372,391)(372,287)(382,287){5}
wire [7:0] w65;    //: /sn:0 {0}(#:227,344)(227,399){1}
//: {2}(229,401)(#:2132,401){3}
//: {4}(225,401)(122,401)(122,321)(132,321){5}
wire [7:0] w56;    //: /sn:0 {0}(#:472,748)(472,801){1}
//: {2}(474,803)(#:1543,803)(1543,435)(#:2132,435){3}
//: {4}(470,803)(373,803)(373,686)(383,686){5}
wire [7:0] w3;    //: /sn:0 {0}(#:481,19)(481,78){1}
wire [7:0] w0;    //: /sn:0 {0}(#:472,551)(472,606){1}
//: {2}(474,608)(1582,608)(1582,421)(#:2132,421){3}
//: {4}(#:470,608)(372,608)(372,494)(382,494){5}
wire [7:0] w22;    //: /sn:0 {0}(#:226,92)(#:226,146){1}
wire w42;    //: /sn:0 {0}(-228,-134)(-26,-134)(-26,249)(398,249)(398,254){1}
wire [7:0] w18;    //: /sn:0 {0}(#:227,551)(227,615){1}
//: {2}(229,617)(#:1567,617)(1567,415)(#:2132,415){3}
//: {4}(225,617)(109,617)(109,529)(119,529){5}
wire w23;    //: /sn:0 {0}(-188,87)(-188,-101)(-228,-101){1}
wire [7:0] w84;    //: /sn:0 {0}(#:412,676)(472,676)(#:472,727){1}
wire [7:0] w21;    //: /sn:0 {0}(#:471,107)(#:471,146){1}
wire [7:0] w24;    //: /sn:0 {0}(#:411,277)(472,277)(#:472,323){1}
wire [7:0] w1;    //: /sn:0 {0}(#:227,748)(227,811){1}
//: {2}(229,813)(#:1532,813)(1532,428)(#:2132,428){3}
//: {4}(225,813)(#:112,813)(112,727)(122,727){5}
wire [7:0] w46;    //: /sn:0 {0}(236,63)(#:236,12){1}
wire w17;    //: /sn:0 {0}(-228,-141)(-58,-141)(-58,273)(148,273)(148,288){1}
wire [7:0] w80;    //: /sn:0 {0}(#:151,717)(227,717)(#:227,727){1}
wire w48;    //: /sn:0 {0}(203,79)(115,79)(115,53){1}
wire w11;    //: /sn:0 {0}(185,-1)(213,-1){1}
wire w41;    //: /sn:0 {0}(135,496)(135,484)(-114,484)(-114,-128)(-228,-128){1}
wire w47;    //: /sn:0 {0}(-228,-114)(-179,-114)(-179,679)(138,679)(138,694){1}
wire w83;    //: /sn:0 {0}(-228,-108)(-142,-108)(-142,638)(399,638)(399,653){1}
wire [7:0] w15;    //: /sn:0 {0}(#:1673,441)(2132,441){1}
wire [7:0] w5;    //: /sn:0 {0}(#:227,323)(227,311)(#:161,311){1}
wire w38;    //: /sn:0 {0}(398,461)(398,457)(-88,457)(-88,-121)(-228,-121){1}
wire [7:0] w76;    //: /sn:0 {0}(#:411,484)(472,484)(#:472,530){1}
wire w26;    //: /sn:0 {0}(113,32)(113,-94)(-228,-94){1}
wire [7:0] w40;    //: /sn:0 {0}(#:227,530)(227,519)(#:148,519){1}
//: enddecls

  //: joint g75 (Clock) @(171, 333) /w:[ 20 22 -1 19 ]
  //: joint g44 (Register_input) @(23, 707) /w:[ 26 28 25 -1 ]
  //: IN g116 (Accumulator_input) @(226,-403) /sn:0 /R:3 /w:[ 1 ]
  //: GROUND g4 (w55) @(291,338) /sn:0 /R:1 /w:[ 0 ]
  //: GROUND g8 (w60) @(295,742) /sn:0 /R:1 /w:[ 0 ]
  //: joint g47 (w18) @(227, 617) /w:[ 2 1 4 -1 ]
  _GGREG8 #(10, 10, 20) B (.Q(w65), .D(w5), .EN(w55), .CLR(_CLR), .CK(Clock));   //: @(227,333) /w:[ 0 0 1 13 21 ]
  //: GROUND g3 (w54) @(546,161) /sn:0 /R:1 /w:[ 0 ]
  _GGOR2 #(6) g90 (.I0(Accumulator_input_choose), .I1(w26), .Z(w48));   //: @(115,43) /sn:0 /R:3 /w:[ 0 0 1 ]
  //: GROUND g2 (w52) @(287,161) /sn:0 /R:1 /w:[ 0 ]
  //: joint g74 (Clock) @(171, 156) /w:[ 24 -1 26 23 ]
  //: joint g23 (_CLR) @(337, 535) /w:[ -1 15 16 18 ]
  _GGREG8 #(10, 10, 20) F (.Q(Flag_output), .D(w21), .EN(w54), .CLR(_CLR), .CK(Clock));   //: @(471,156) /w:[ 3 1 1 0 11 ]
  //: joint g77 (Clock) @(425, 540) /w:[ 14 13 -1 16 ]
  //: joint g39 (Register_input) @(44, 301) /w:[ 1 2 4 -1 ]
  //: joint g24 (_CLR) @(337, 328) /w:[ -1 11 12 14 ]
  //: IN g86 (Flag_input_choose) @(480,-653) /sn:0 /R:3 /w:[ 0 ]
  _GGMUX2x8 #(8, 8) g60 (.I0(w56), .I1(Register_input), .S(w83), .Z(w84));   //: @(399,676) /sn:0 /R:1 /w:[ 5 29 1 0 ] /ss:1 /do:0
  _GGREG8 #(10, 10, 20) A (.Q(Accumulator_output), .D(w22), .EN(w52), .CLR(_CLR), .CK(Clock));   //: @(226,156) /w:[ 9 1 1 9 25 ]
  _GGMUX2x8 #(8, 8) g82 (.I0(Flag_output), .I1(w3), .S(Flag_input_choose), .Z(w21));   //: @(471,94) /sn:0 /w:[ 5 1 5 0 ] /ss:0 /do:0
  //: IN g70 (Clock) @(-99,-266) /sn:0 /w:[ 27 ]
  //: IN g18 (_CLR) @(-66,-300) /sn:0 /w:[ 5 ]
  //: joint g65 (w56) @(472, 803) /w:[ 2 1 4 -1 ]
  //: joint g64 (w13) @(472, 391) /w:[ 2 1 4 -1 ]
  _GGMUX2x8 #(8, 8) g49 (.I0(Accumulator_output), .I1(w46), .S(w48), .Z(w22));   //: @(226,79) /sn:0 /w:[ 0 0 0 0 ] /ss:0 /do:0
  //: OUT g50 (Register_output1) @(2512,425) /sn:0 /w:[ 1 ]
  //: GROUND g6 (w58) @(286,545) /sn:0 /R:1 /w:[ 0 ]
  //: joint g68 (Register_input) @(-52, 509) /w:[ 20 22 19 -1 ]
  _GGMUX2x8 #(8, 8) g58 (.I0(w0), .I1(Register_input), .S(w38), .Z(w76));   //: @(398,484) /sn:0 /R:1 /w:[ 5 23 0 0 ] /ss:1 /do:0
  _GGMUX2x8 #(8, 8) g56 (.I0(w18), .I1(Register_input), .S(w41), .Z(w40));   //: @(135,519) /sn:0 /R:1 /w:[ 5 21 0 1 ] /ss:1 /do:0
  //: IN g73 (Register_input_choose) @(-503,-118) /sn:0 /w:[ 0 ]
  //: joint g35 (Register_input) @(-340, -52) /w:[ 8 -1 14 7 ]
  //: GROUND g7 (w59) @(524,545) /sn:0 /R:1 /w:[ 0 ]
  //: GROUND g9 (w61) @(531,742) /sn:0 /R:1 /w:[ 0 ]
  _GGMUX2x8 #(8, 8) g59 (.I0(w1), .I1(Register_input), .S(w47), .Z(w80));   //: @(138,717) /sn:0 /R:1 /w:[ 5 27 1 0 ] /ss:1 /do:0
  //: joint g22 (_CLR) @(337, 151) /w:[ -1 7 8 10 ]
  //: IN g71 (Register_output_choose1) @(2084,-150) /sn:0 /w:[ 0 ]
  //: joint g31 (_CLR) @(337, -300) /w:[ 3 -1 4 6 ]
  //: joint g67 (w0) @(472, 608) /w:[ 2 1 4 -1 ]
  //: joint g83 (Flag_input_choose) @(421, 6) /w:[ 2 1 -1 4 ]
  //: joint g41 (Accumulator_input_choose) @(118, 1) /w:[ 2 4 -1 1 ]
  //: joint g45 (Register_input_dec) @(-244, -216) /w:[ 2 -1 1 4 ]
  //: IN g36 (Register_input_dec) @(-503,-216) /sn:0 /w:[ 0 ]
  //: joint g81 (Clock) @(425, 425) /w:[ -1 6 5 12 ]
  //: joint g69 (Accumulator_output) @(226, 217) /w:[ 2 8 1 -1 ]
  //: joint g42 (Register_input) @(-340, 301) /w:[ 5 6 -1 16 ]
  _GGAND2 #(6) g40 (.I0(!Register_input_dec), .I1(Accumulator_input_choose), .Z(w11));   //: @(175,-1) /sn:0 /w:[ 3 3 0 ]
  _GGDECODER8 #(6, 6) g52 (.I(Register_input_choose), .E(Register_input_dec), .Z0(w17), .Z1(w42), .Z2(w41), .Z3(w38), .Z4(w47), .Z5(w83), .Z6(w23), .Z7(w26));   //: @(-244,-118) /sn:0 /R:1 /w:[ 1 5 0 0 1 1 0 0 1 1 ] /ss:1 /do:1
  //: joint g66 (w1) @(227, 813) /w:[ 2 1 4 -1 ]
  _GGMUX2x8 #(8, 8) g46 (.I0(w65), .I1(Register_input), .S(w17), .Z(w5));   //: @(148,311) /sn:0 /R:1 /w:[ 5 0 1 1 ] /ss:1 /do:0
  //: IN g34 (Register_input) @(-503,-52) /sn:0 /w:[ 15 ]
  //: joint g57 (Accumulator_output) @(320, 217) /w:[ 4 6 3 -1 ]
  //: joint g84 (Clock) @(425, 333) /w:[ 8 10 -1 7 ]
  //: OUT g118 (Accumulator_output) @(320,-653) /sn:0 /R:1 /w:[ 7 ]
  //: GROUND g5 (w57) @(540,338) /sn:0 /R:1 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) H (.Q(w1), .D(w80), .EN(w60), .CLR(_CLR), .CK(Clock));   //: @(227,737) /w:[ 0 1 1 19 29 ]
  _GGMUX8x8 #(20, 20) g61 (.I0(w65), .I1(w13), .I2(w18), .I3(w0), .I4(w1), .I5(w56), .I6(w15), .I7(Accumulator_output), .S(Register_output_choose1), .Z(Register_output1));   //: @(2148,425) /sn:0 /R:1 /w:[ 3 3 3 3 3 3 1 5 1 0 ] /ss:1 /do:1
  //: joint g21 (_CLR) @(560, 151) /w:[ -1 2 1 20 ]
  //: joint g19 (_CLR) @(560, 535) /w:[ -1 25 26 28 ]
  _GGREG8 #(10, 10, 20) D (.Q(w18), .D(w40), .EN(w58), .CLR(_CLR), .CK(Clock));   //: @(227,540) /w:[ 0 0 1 17 0 ]
  _GGREG8 #(10, 10, 20) C (.Q(w13), .D(w24), .EN(w57), .CLR(_CLR), .CK(Clock));   //: @(472,333) /w:[ 0 1 1 23 9 ]
  //: joint g79 (Clock) @(171, 425) /w:[ 4 18 -1 3 ]
  //: joint g20 (_CLR) @(560, 328) /w:[ -1 21 22 24 ]
  //: joint g115 (Register_input) @(246, -52) /w:[ 10 -1 9 12 ]
  //: OUT g78 (Flag_output) @(655,-648) /sn:0 /R:1 /w:[ 0 ]
  //: joint g43 (Register_input) @(-340, 509) /w:[ 18 17 -1 24 ]
  //: frame g0 @(150,111) /sn:0 /wi:399 /ht:676 /tx:"Main registers"
  _GGMUX2x8 #(8, 8) g38 (.I0(Register_input), .I1(Accumulator_input), .S(w11), .Z(w46));   //: @(236,-1) /sn:0 /w:[ 13 0 1 1 ] /ss:0 /do:1
  _GGMUX2x8 #(8, 8) g48 (.I0(w13), .I1(Register_input), .S(w42), .Z(w24));   //: @(398,277) /sn:0 /R:1 /w:[ 5 3 1 0 ] /ss:1 /do:0
  _GGREG8 #(10, 10, 20) E (.Q(w0), .D(w76), .EN(w59), .CLR(_CLR), .CK(Clock));   //: @(472,540) /w:[ 0 1 1 27 15 ]
  //: joint g62 (w65) @(227, 401) /w:[ 2 1 4 -1 ]
  _GGMUX2x8 #(8, 8) g37 (.I0(Register_input), .I1(Flag_input), .S(Flag_input_choose), .Z(w3));   //: @(481,6) /sn:0 /w:[ 11 0 3 0 ] /ss:0 /do:1
  //: joint g55 (Flag_output) @(471, 204) /w:[ 1 2 4 -1 ]
  _GGREG8 #(10, 10, 20) L (.Q(w56), .D(w84), .EN(w61), .CLR(_CLR), .CK(Clock));   //: @(472,737) /w:[ 0 1 1 29 17 ]
  //: IN g88 (Accumulator_input_choose) @(118,-653) /sn:0 /R:3 /w:[ 5 ]
  //: IN g80 (Flag_input) @(567,-490) /sn:0 /R:3 /w:[ 1 ]
  //: joint g76 (Clock) @(171, 540) /w:[ 1 2 -1 28 ]

endmodule
//: /netlistEnd

//: /netlistBegin make_negative
module make_negative(Output0, Input0);
//: interface  /sz:(101, 47) /bd:[ Ti0>Input0[7:0](21/101) Bo0<Output0[7:0](21/101) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply0 w0;    //: /sn:0 {0}(469,241)(417,241)(417,223){1}
//: {2}(419,221)(434,221){3}
//: {4}(438,221)(469,221){5}
//: {6}(436,223)(436,231)(469,231){7}
//: {8}(415,221)(398,221){9}
//: {10}(396,219)(396,193){11}
//: {12}(398,191)(418,191){13}
//: {14}(422,191)(449,191){15}
//: {16}(453,191)(469,191){17}
//: {18}(451,193)(451,201)(469,201){19}
//: {20}(420,193)(420,211)(469,211){21}
//: {22}(394,191)(284,191){23}
//: {24}(396,223)(396,251)(469,251){25}
output [7:0] Output0;    //: /sn:0 {0}(#:566,168)(819,168){1}
input [7:0] Input0;    //: /sn:0 {0}(537,152)(#:428,152){1}
supply0 w1;    //: /sn:0 {0}(551,113)(551,144){1}
supply1 w2;    //: /sn:0 {0}(212,152)(212,261)(469,261){1}
wire w16;    //: /sn:0 {0}(611,203)(551,203)(551,192){1}
wire [7:0] w5;    //: /sn:0 {0}(#:475,226)(522,226)(522,184)(537,184){1}
//: enddecls

  //: joint g8 (w0) @(451, 191) /w:[ 16 -1 15 18 ]
  //: VDD g4 (w2) @(223,152) /sn:0 /w:[ 0 ]
  //: GROUND g3 (w1) @(551,107) /sn:0 /R:2 /w:[ 0 ]
  //: GROUND g2 (w0) @(278,191) /sn:0 /R:3 /w:[ 23 ]
  //: OUT g1 (Output0) @(816,168) /sn:0 /w:[ 1 ]
  //: joint g10 (w0) @(396, 191) /w:[ 12 -1 22 11 ]
  _GGADD8 #(68, 70, 62, 64) g6 (.A(w5), .B(Input0), .S(Output0), .CI(w1), .CO(w16));   //: @(553,168) /sn:0 /R:1 /w:[ 1 0 0 1 1 ]
  //: joint g9 (w0) @(420, 191) /w:[ 14 -1 13 20 ]
  //: LED g7 (w16) @(618,203) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g12 (w0) @(417, 221) /w:[ 2 -1 8 1 ]
  //: joint g11 (w0) @(436, 221) /w:[ 4 -1 3 6 ]
  assign w5 = {w0, w0, w0, w0, w0, w0, w0, w2}; //: CONCAT g5  @(474,226) /sn:0 /w:[ 0 17 19 21 5 7 0 25 1 ] /dr:0 /tp:0 /drp:1
  //: IN g0 (Input0) @(426,152) /sn:0 /w:[ 1 ]
  //: joint g13 (w0) @(396, 221) /w:[ 9 10 -1 24 ]

endmodule
//: /netlistEnd

//: /netlistBegin set_flags
module set_flags(x6_zero_flag, x2_parity_overflow_flag, x2_input_01, x1_subtract_flag_set, x2_set_01, x1_subtract_flag, x6_set_01, x6_set_by_bits, x0_carry_flag_set, x4_set_01, x7_sign_flag, x4_input_01, x4_set_by_bits, x4_halfcarry_flag, x6_zero_flag_set, x4_halfcarry_flag_set, x0_input_01, x6_input_by_bits, x1_input_01, x2_set_overflow, x0_input_by_bits, x2_input_parity, x2_input_overflow, x7_input_01, x7_set_01, x7_sign_flag_set, x2_parity_overflow_flag_set, x6_input_01, x1_set_01, x7_set_by_bits, x0_carry_flag, x0_set_by_bits, x4_input_by_bits, x0_set_01, x2_set_parity, x7_input_by_bits);
//: interface  /sz:(393, 400) /bd:[ Li0>x7_set_by_bits(384/400) Li1>x7_set_01(368/400) Li2>x7_input_by_bits[7:0](352/400) Li3>x7_input_01(336/400) Li4>x6_set_by_bits(320/400) Li5>x6_set_01(304/400) Li6>x6_input_by_bits[7:0](288/400) Li7>x6_input_01(272/400) Li8>x4_set_by_bits(256/400) Li9>x4_set_01(240/400) Li10>x4_input_by_bits(224/400) Li11>x4_input_01(208/400) Li12>x2_set_parity(192/400) Li13>x2_set_overflow(176/400) Li14>x2_set_01(160/400) Li15>x2_input_parity[7:0](144/400) Li16>x2_input_overflow(128/400) Li17>x2_input_01(112/400) Li18>x1_set_01(96/400) Li19>x1_input_01(80/400) Li20>x0_set_by_bits(64/400) Li21>x0_set_01(48/400) Li22>x0_input_by_bits(32/400) Li23>x0_input_01(16/400) Ro0<x7_sign_flag_set(192/400) Ro1<x7_sign_flag(176/400) Ro2<x6_zero_flag_set(160/400) Ro3<x6_zero_flag(144/400) Ro4<x4_halfcarry_flag_set(128/400) Ro5<x4_halfcarry_flag(112/400) Ro6<x2_parity_overflow_flag_set(96/400) Ro7<x2_parity_overflow_flag(80/400) Ro8<x1_subtract_flag_set(64/400) Ro9<x1_subtract_flag(48/400) Ro10<x0_carry_flag_set(32/400) Ro11<x0_carry_flag(16/400) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output x1_subtract_flag;    //: /sn:0 {0}(197,113)(938,113)(938,113)(991,113){1}
input [7:0] x2_input_parity;    //: /sn:0 {0}(#:195,290)(175,290)(175,255)(128,255){1}
input x0_input_01;    //: /sn:0 {0}(105,-57)(168,-57)(168,-57)(183,-57){1}
input x2_set_01;    //: /sn:0 {0}(128,363)(334,363){1}
//: {2}(338,363)(375,363){3}
//: {4}(336,365)(336,381)(410,381){5}
input x7_input_01;    //: /sn:0 {0}(397,736)(310,736)(310,736)(196,736){1}
input x0_input_by_bits;    //: /sn:0 {0}(183,-37)(120,-37)(120,-37)(105,-37){1}
input x4_set_by_bits;    //: /sn:0 {0}(126,520)(183,520){1}
//: {2}(187,520)(207,520){3}
//: {4}(185,522)(185,550)(207,550){5}
output x0_carry_flag;    //: /sn:0 {0}(212,-47)(234,-47)(234,7)(991,7){1}
output x7_sign_flag;    //: /sn:0 {0}(426,746)(1075,746)(1075,746)(991,746){1}
output x0_carry_flag_set;    //: /sn:0 {0}(172,27)(204,27)(204,27)(991,27){1}
output x6_zero_flag;    //: /sn:0 {0}(991,634)(366,634)(366,634)(351,634){1}
input x4_input_01;    //: /sn:0 {0}(124,489)(239,489){1}
input x2_set_overflow;    //: /sn:0 {0}(410,391)(395,391)(395,406){1}
//: {2}(397,408)(547,408)(547,254){3}
//: {4}(393,408)(128,408){5}
output x4_halfcarry_flag_set;    //: /sn:0 {0}(993,553)(878,553)(878,553)(228,553){1}
input x6_set_by_bits;    //: /sn:0 {0}(163,694)(184,694){1}
//: {2}(188,694)(259,694){3}
//: {4}(186,692)(186,675)(259,675){5}
output x7_sign_flag_set;    //: /sn:0 {0}(377,810)(434,810)(434,766)(991,766){1}
output x1_subtract_flag_set;    //: /sn:0 {0}(197,133)(481,133)(481,133)(991,133){1}
input x1_set_01;    //: /sn:0 {0}(129,133)(127,133)(127,133)(176,133){1}
input [7:0] x7_input_by_bits;    //: /sn:0 {0}(#:196,756)(223,756){1}
//: {2}(224,756)(#:235,756){3}
input x2_set_parity;    //: /sn:0 {0}(128,386)(295,386){1}
//: {2}(299,386)(410,386){3}
//: {4}(297,384)(297,368)(375,368){5}
output x2_parity_overflow_flag;    //: /sn:0 {0}(560,231)(596,231)(596,241)(991,241){1}
input x2_input_01;    //: /sn:0 {0}(427,231)(128,231){1}
input x4_set_01;    //: /sn:0 {0}(127,555)(174,555){1}
//: {2}(178,555)(193,555)(193,555)(207,555){3}
//: {4}(176,553)(176,525)(207,525){5}
output x6_zero_flag_set;    //: /sn:0 {0}(280,692)(369,692)(369,654)(991,654){1}
input x0_set_01;    //: /sn:0 {0}(151,-6)(131,-6){1}
//: {2}(127,-6)(105,-6){3}
//: {4}(129,-4)(129,24)(151,24){5}
input x2_input_overflow;    //: /sn:0 {0}(128,209)(515,209)(515,221)(531,221){1}
input x7_set_by_bits;    //: /sn:0 {0}(355,791)(310,791)(310,810){1}
//: {2}(312,812)(356,812){3}
//: {4}(308,812)(301,812)(301,812)(196,812){5}
output x4_halfcarry_flag;    //: /sn:0 {0}(993,533)(290,533)(290,479)(268,479){1}
output x2_parity_overflow_flag_set;    //: /sn:0 {0}(431,386)(596,386)(596,261)(991,261){1}
input x4_input_by_bits;    //: /sn:0 {0}(129,469)(239,469){1}
input x1_input_01;    //: /sn:0 {0}(176,113)(135,113)(135,113)(129,113){1}
input x7_set_01;    //: /sn:0 {0}(196,786)(312,786)(312,786)(330,786){1}
//: {2}(334,786)(355,786){3}
//: {4}(332,788)(332,807)(356,807){5}
input [7:0] x6_input_by_bits;    //: /sn:0 {0}(211,644)(#:163,644){1}
input x6_set_01;    //: /sn:0 {0}(259,670)(222,670){1}
//: {2}(218,670)(163,670){3}
//: {4}(220,672)(220,689)(259,689){5}
input x6_input_01;    //: /sn:0 {0}(163,624)(213,624)(213,624)(322,624){1}
input x0_set_by_bits;    //: /sn:0 {0}(151,29)(137,29)(137,29)(122,29){1}
//: {2}(120,27)(120,-1)(151,-1){3}
//: {4}(118,29)(105,29){5}
wire w16;    //: /sn:0 {0}(297,258)(279,258)(279,258)(259,258){1}
wire w13;    //: /sn:0 {0}(238,315)(219,315)(219,315)(201,315){1}
wire w6;    //: /sn:0 {0}(232,644)(307,644)(307,644)(322,644){1}
wire w7;    //: /sn:0 {0}(238,260)(217,260)(217,265)(201,265){1}
wire w25;    //: /sn:0 {0}(297,303)(271,303)(271,318)(259,318){1}
wire w4;    //: /sn:0 {0}(172,-3)(199,-3)(199,-24){1}
wire w22;    //: /sn:0 {0}(297,298)(276,298)(276,298)(259,298){1}
wire w0;    //: /sn:0 {0}(360,264)(387,264)(387,251)(427,251){1}
wire w3;    //: /sn:0 {0}(280,673)(338,673)(338,657){1}
wire w18;    //: /sn:0 {0}(456,241)(531,241){1}
wire w19;    //: /sn:0 {0}(297,263)(276,263)(276,278)(259,278){1}
wire w12;    //: /sn:0 {0}(238,300)(212,300)(212,305)(201,305){1}
wire w10;    //: /sn:0 {0}(238,280)(215,280)(215,285)(201,285){1}
wire w21;    //: /sn:0 {0}(339,266)(324,266)(324,301)(318,301){1}
wire w1;    //: /sn:0 {0}(238,255)(220,255)(220,255)(201,255){1}
wire w8;    //: /sn:0 {0}(397,756)(310,756)(310,744)(224,744)(224,751){1}
wire w17;    //: /sn:0 {0}(339,261)(318,261){1}
wire w14;    //: /sn:0 {0}(238,320)(215,320)(215,325)(201,325){1}
wire w11;    //: /sn:0 {0}(238,295)(218,295)(218,295)(201,295){1}
wire w2;    //: /sn:0 {0}(413,769)(413,789)(376,789){1}
wire w15;    //: /sn:0 {0}(228,523)(255,523)(255,502){1}
wire w5;    //: /sn:0 {0}(396,366)(443,366)(443,264){1}
wire w9;    //: /sn:0 {0}(238,275)(219,275)(219,275)(201,275){1}
//: enddecls

  //: OUT g8 (x6_zero_flag) @(988,634) /sn:0 /w:[ 0 ]
  //: OUT g4 (x2_parity_overflow_flag) @(988,241) /sn:0 /w:[ 1 ]
  //: IN g44 (x2_input_01) @(126,231) /sn:0 /w:[ 1 ]
  _GGMUX2 #(8, 8) g16 (.I0(w8), .I1(x7_input_01), .S(w2), .Z(x7_sign_flag));   //: @(413,746) /sn:0 /R:1 /w:[ 0 0 0 0 ] /ss:0 /do:0
  //: OUT g3 (x1_subtract_flag_set) @(988,133) /sn:0 /w:[ 1 ]
  //: IN g47 (x2_set_01) @(126,363) /sn:0 /w:[ 0 ]
  _GGNOR1x8 #(1) g26 (.I0(x6_input_by_bits), .Z(w6));   //: @(222,644) /sn:0 /w:[ 0 0 ]
  _GGAND2 #(6) g17 (.I0(x7_set_01), .I1(!x7_set_by_bits), .Z(w2));   //: @(366,789) /sn:0 /w:[ 3 0 1 ]
  //: OUT g2 (x1_subtract_flag) @(988,113) /sn:0 /w:[ 1 ]
  //: joint g74 (x4_set_01) @(176, 555) /w:[ 2 4 1 -1 ]
  //: IN g23 (x6_set_01) @(161,670) /sn:0 /w:[ 3 ]
  //: joint g30 (x6_set_01) @(220, 670) /w:[ 1 -1 2 4 ]
  //: IN g24 (x6_set_by_bits) @(161,694) /sn:0 /w:[ 0 ]
  //: OUT g1 (x0_carry_flag_set) @(988,27) /sn:0 /w:[ 1 ]
  _GGMUX2 #(8, 8) g39 (.I0(x0_input_by_bits), .I1(x0_input_01), .S(w4), .Z(x0_carry_flag));   //: @(199,-47) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:0
  _GGNXOR2 #(6) g60 (.I0(w17), .I1(w21), .Z(w0));   //: @(350,264) /sn:0 /w:[ 0 0 0 ]
  //: joint g29 (x6_set_by_bits) @(186, 694) /w:[ 2 4 1 -1 ]
  //: IN g51 (x4_set_01) @(125,555) /sn:0 /w:[ 0 ]
  _GGMUX2 #(8, 8) g70 (.I0(x4_input_01), .I1(x4_input_by_bits), .S(w15), .Z(x4_halfcarry_flag));   //: @(255,479) /sn:0 /R:1 /w:[ 1 1 1 1 ] /ss:0 /do:0
  _GGOR2 #(6) g18 (.I0(x7_set_01), .I1(x7_set_by_bits), .Z(x7_sign_flag_set));   //: @(367,810) /sn:0 /w:[ 5 3 0 ]
  _GGMUX2 #(8, 8) g25 (.I0(w6), .I1(x6_input_01), .S(w3), .Z(x6_zero_flag));   //: @(338,634) /sn:0 /R:1 /w:[ 1 1 1 1 ] /ss:0 /do:0
  //: OUT g10 (x7_sign_flag) @(988,746) /sn:0 /w:[ 1 ]
  assign w8 = x7_input_by_bits[7]; //: TAP g65 @(224,754) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:0
  //: joint g64 (x2_set_parity) @(297, 386) /w:[ 2 4 1 -1 ]
  //: IN g49 (x4_input_01) @(122,489) /sn:0 /w:[ 0 ]
  //: joint g72 (x4_set_by_bits) @(185, 520) /w:[ 2 -1 1 4 ]
  //: IN g50 (x4_set_by_bits) @(124,520) /sn:0 /w:[ 0 ]
  //: OUT g6 (x4_halfcarry_flag) @(990,533) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g73 (.I0(x4_set_by_bits), .I1(!x4_set_01), .Z(w15));   //: @(218,523) /sn:0 /w:[ 3 5 0 ]
  _GGMUX2 #(8, 8) g68 (.I0(w18), .I1(x2_input_overflow), .S(x2_set_overflow), .Z(x2_parity_overflow_flag));   //: @(547,231) /sn:0 /R:1 /w:[ 1 1 3 0 ] /ss:0 /do:0
  _GGXOR2 #(8) g58 (.I0(w16), .I1(w19), .Z(w17));   //: @(308,261) /sn:0 /w:[ 0 0 1 ]
  _GGXOR2 #(8) g56 (.I0(w11), .I1(w12), .Z(w22));   //: @(249,298) /sn:0 /w:[ 0 0 1 ]
  //: OUT g9 (x6_zero_flag_set) @(988,654) /sn:0 /w:[ 1 ]
  //: OUT g7 (x4_halfcarry_flag_set) @(990,553) /sn:0 /w:[ 0 ]
  //: IN g35 (x0_input_01) @(103,-57) /sn:0 /w:[ 0 ]
  _GGOR2 #(6) g71 (.I0(x4_set_by_bits), .I1(x4_set_01), .Z(x4_halfcarry_flag_set));   //: @(218,553) /sn:0 /w:[ 5 3 1 ]
  _GGXOR2 #(8) g59 (.I0(w22), .I1(w25), .Z(w21));   //: @(308,301) /sn:0 /w:[ 0 0 1 ]
  //: IN g22 (x6_input_by_bits) @(161,644) /sn:0 /w:[ 1 ]
  //: IN g31 (x1_input_01) @(127,113) /sn:0 /w:[ 1 ]
  //: IN g67 (x2_set_overflow) @(126,408) /sn:0 /w:[ 5 ]
  _GGXOR2 #(8) g54 (.I0(w1), .I1(w7), .Z(w16));   //: @(249,258) /sn:0 /w:[ 0 0 1 ]
  _GGMUX2 #(8, 8) g45 (.I0(w0), .I1(x2_input_01), .S(w5), .Z(w18));   //: @(443,241) /sn:0 /R:1 /w:[ 1 0 1 0 ] /ss:0 /do:0
  _GGOR1 #(1) g33 (.I0(x1_set_01), .Z(x1_subtract_flag_set));   //: @(187,133) /sn:0 /w:[ 1 0 ]
  //: IN g36 (x0_input_by_bits) @(103,-37) /sn:0 /w:[ 1 ]
  _GGOR2 #(6) g41 (.I0(x0_set_01), .I1(x0_set_by_bits), .Z(x0_carry_flag_set));   //: @(162,27) /sn:0 /w:[ 5 0 0 ]
  //: joint g69 (x2_set_overflow) @(395, 408) /w:[ 2 1 4 -1 ]
  //: IN g52 (x2_input_parity) @(126,255) /sn:0 /w:[ 1 ]
  _GGAND2 #(6) g40 (.I0(x0_set_01), .I1(!x0_set_by_bits), .Z(w4));   //: @(162,-3) /sn:0 /w:[ 0 3 0 ]
  //: joint g42 (x0_set_01) @(129, -6) /w:[ 1 -1 2 4 ]
  //: IN g66 (x2_input_overflow) @(126,209) /sn:0 /w:[ 0 ]
  //: IN g12 (x7_input_01) @(194,736) /sn:0 /w:[ 1 ]
  _GGXOR2 #(8) g57 (.I0(w13), .I1(w14), .Z(w25));   //: @(249,318) /sn:0 /w:[ 0 0 1 ]
  assign {w14, w13, w12, w11, w10, w9, w7, w1} = x2_input_parity; //: CONCAT g46  @(196,290) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  _GGOR2 #(6) g28 (.I0(x6_set_01), .I1(x6_set_by_bits), .Z(x6_zero_flag_set));   //: @(270,692) /sn:0 /w:[ 5 3 0 ]
  _GGOR1 #(1) g34 (.I0(x1_input_01), .Z(x1_subtract_flag));   //: @(187,113) /sn:0 /w:[ 0 0 ]
  //: IN g14 (x7_set_01) @(194,786) /sn:0 /w:[ 0 ]
  //: OUT g11 (x7_sign_flag_set) @(988,766) /sn:0 /w:[ 1 ]
  //: OUT g5 (x2_parity_overflow_flag_set) @(988,261) /sn:0 /w:[ 1 ]
  _GGAND2 #(6) g61 (.I0(x2_set_01), .I1(!x2_set_parity), .Z(w5));   //: @(386,366) /sn:0 /w:[ 3 5 0 ]
  //: IN g21 (x6_input_01) @(161,624) /sn:0 /w:[ 0 ]
  //: joint g19 (x7_set_by_bits) @(310, 812) /w:[ 2 1 4 -1 ]
  //: joint g20 (x7_set_01) @(332, 786) /w:[ 2 -1 1 4 ]
  //: IN g32 (x1_set_01) @(127,133) /sn:0 /w:[ 0 ]
  //: joint g63 (x2_set_01) @(336, 363) /w:[ 2 -1 1 4 ]
  //: IN g15 (x7_set_by_bits) @(194,812) /sn:0 /w:[ 5 ]
  //: OUT g0 (x0_carry_flag) @(988,7) /sn:0 /w:[ 1 ]
  //: IN g38 (x0_set_by_bits) @(103,29) /sn:0 /w:[ 5 ]
  //: joint g43 (x0_set_by_bits) @(120, 29) /w:[ 1 2 4 -1 ]
  _GGAND2 #(6) g27 (.I0(x6_set_01), .I1(!x6_set_by_bits), .Z(w3));   //: @(270,673) /sn:0 /w:[ 0 5 0 ]
  //: IN g48 (x4_input_by_bits) @(127,469) /sn:0 /w:[ 0 ]
  _GGOR3 #(8) g62 (.I0(x2_set_01), .I1(x2_set_parity), .I2(x2_set_overflow), .Z(x2_parity_overflow_flag_set));   //: @(421,386) /sn:0 /w:[ 5 3 0 0 ]
  //: IN g37 (x0_set_01) @(103,-6) /sn:0 /w:[ 3 ]
  _GGXOR2 #(8) g55 (.I0(w9), .I1(w10), .Z(w19));   //: @(249,278) /sn:0 /w:[ 0 0 1 ]
  //: IN g53 (x2_set_parity) @(126,386) /sn:0 /w:[ 0 ]
  //: IN g13 (x7_input_by_bits) @(194,756) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin registers_old
module registers_old(Accumulator_input, Register_output2, Register_output_choose2, Flag_output, Flag_input, Flag_input_choose, Register_reset, Register_output1, Register_input_choose, Register_output_choose1, Register_input, Accumulator_output, Use_shadow_reg, Accumulator_input_choose);
//: interface  /sz:(441, 192) /bd:[ Li0>Use_shadow_reg(160/192) Li1>Register_reset(144/192) Li2>Register_output_choose2[7:0](128/192) Li3>Register_output_choose1[7:0](112/192) Li4>Register_input_choose[7:0](96/192) Li5>Register_input[7:0](80/192) Li6>Flag_input_choose(64/192) Li7>Flag_input[7:0](48/192) Li8>Accumulator_input_choose(32/192) Li9>Accumulator_input[7:0](16/192) Ro0<Register_output2[7:0](64/192) Ro1<Register_output1[7:0](48/192) Ro2<Flag_output[7:0](32/192) Ro3<Accumulator_output[7:0](16/192) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] Register_output_choose2;    //: /sn:0 {0}(#:1632,-198)(1739,-198){1}
//: {2}(1740,-198)(1770,-198){3}
//: {4}(1771,-198)(1787,-198){5}
input [7:0] Register_input;    //: /sn:0 {0}(#:-386,-52)(-342,-52){1}
//: {2}(-338,-52)(234,-52){3}
//: {4}(238,-52)(453,-52){5}
//: {6}(457,-52)(998,-52){7}
//: {8}(1002,-52)(1220,-52)(#:1220,-10){9}
//: {10}(1000,-50)(1000,-16){11}
//: {12}(455,-50)(455,-10){13}
//: {14}(236,-50)(236,-17){15}
//: {16}(-340,-50)(-340,309){17}
//: {18}(-338,311)(225,311){19}
//: {20}(229,311)(444,311){21}
//: {22}(448,311)(989,311){23}
//: {24}(#:993,311)(1210,311)(1210,323){25}
//: {26}(991,313)(#:991,323){27}
//: {28}(446,313)(#:446,323){29}
//: {30}(227,313)(#:227,323){31}
//: {32}(#:-340,313)(-340,516){33}
//: {34}(-338,518)(225,518){35}
//: {36}(#:229,518)(444,518){37}
//: {38}(#:448,518)(989,518){39}
//: {40}(#:993,518)(1211,518)(1211,530){41}
//: {42}(991,520)(991,530){43}
//: {44}(446,520)(446,530){45}
//: {46}(227,520)(227,530){47}
//: {48}(#:-340,520)(-340,716)(225,716){49}
//: {50}(#:229,716)(444,716){51}
//: {52}(#:448,716)(989,716){53}
//: {54}(#:993,716)(1210,716)(1210,727){55}
//: {56}(991,718)(991,727){57}
//: {58}(446,718)(446,727){59}
//: {60}(227,718)(227,727){61}
input Register_reset;    //: /sn:0 {0}(-49,-300)(-64,-300){1}
output [7:0] Register_output1;    //: /sn:0 {0}(#:2470,61)(#:2817,61){1}
input [7:0] Register_input_choose;    //: /sn:0 {0}(#:-671,-251)(-616,-251){1}
//: {2}(-615,-251)(-549,-251){3}
//: {4}(-548,-251)(-512,-251){5}
output [7:0] Register_output2;    //: /sn:0 {0}(#:2660,255)(2807,255)(2807,254)(2817,254){1}
input Accumulator_input_choose;    //: /sn:0 {0}(197,-649)(197,-512)(242,-512)(242,-497){1}
input [7:0] Flag_input;    //: /sn:0 {0}(#:1200,-10)(1200,-383)(762,-383){1}
//: {2}(760,-385)(#:760,-399){3}
//: {4}(758,-383)(435,-383)(#:435,-10){5}
output [7:0] Accumulator_output;    //: /sn:0 {0}(#:436,-598)(436,-664){1}
output [7:0] Flag_output;    //: /sn:0 {0}(#:1115,-654)(#:1115,-571){1}
input Use_shadow_reg;    //: /sn:0 {0}(264,-484)(272,-484)(272,-492)(656,-492)(656,-556){1}
//: {2}(658,-558)(1092,-558){3}
//: {4}(656,-560)(656,-583){5}
//: {6}(658,-585)(883,-585){7}
//: {8}(656,-587)(656,-622){9}
//: {10}(654,-585)(459,-585){11}
supply0 w80;    //: /sn:0 {0}(265,161)(300,161)(300,336){1}
//: {2}(298,338)(266,338){3}
//: {4}(300,340)(300,543){5}
//: {6}(298,545)(266,545){7}
//: {8}(300,547)(300,740){9}
//: {10}(298,742)(266,742){11}
//: {12}(300,744)(300,854)(611,854){13}
//: {14}(613,852)(613,744){15}
//: {16}(613,740)(613,547){17}
//: {18}(613,543)(613,340){19}
//: {20}(613,336)(613,161)(484,161){21}
//: {22}(611,338)(485,338){23}
//: {24}(611,545)(485,545){25}
//: {26}(611,742)(485,742){27}
//: {28}(613,856)(613,859){29}
//: {30}(615,861)(1064,861){31}
//: {32}(1068,861)(1278,861)(1278,744){33}
//: {34}(1278,740)(1278,547){35}
//: {36}(1278,543)(1278,340){37}
//: {38}(1278,336)(1278,161)(1249,161){39}
//: {40}(1276,338)(1249,338){41}
//: {42}(1276,545)(1250,545){43}
//: {44}(1276,742)(1249,742){45}
//: {46}(1066,859)(1066,744){47}
//: {48}(1066,740)(1066,547){49}
//: {50}(1066,543)(1066,340){51}
//: {52}(1066,336)(1066,161)(1029,161){53}
//: {54}(1064,338)(1030,338){55}
//: {56}(1064,545)(1030,545){57}
//: {58}(1064,742)(1030,742){59}
//: {60}(613,863)(613,925){61}
input [7:0] Register_output_choose1;    //: /sn:0 {0}(#:1578,-150)(1655,-150){1}
//: {2}(1656,-150)(1683,-150){3}
//: {4}(1684,-150)(1699,-150){5}
input [7:0] Accumulator_input;    //: /sn:0 {0}(#:216,-401)(216,-332){1}
//: {2}(#:218,-330)(980,-330)(980,-16){3}
//: {4}(216,-328)(216,-17){5}
input Flag_input_choose;    //: /sn:0 {0}(907,-598)(907,-625){1}
supply1 w40;    //: /sn:0 {0}(-470,-295)(-470,-252){1}
wire [7:0] w16;    //: /sn:0 {0}(#:991,551)(991,569)(1397,569)(1397,41)(1759,41){1}
//: {2}(1763,41)(1801,41){3}
//: {4}(1761,43)(1761,122)(1887,122){5}
wire [7:0] w13;    //: /sn:0 {0}(#:2132,408)(2106,408){1}
//: {2}(2102,408)(1525,408)(#:1525,391)(446,391)(#:446,344){3}
//: {4}(#:2104,410)(2104,514)(2220,514){5}
wire [7:0] w6;    //: /sn:0 {0}(#:1210,344)(1210,351)(1369,351)(1369,34)(1774,34){1}
//: {2}(1778,34)(1801,34){3}
//: {4}(1776,36)(1776,115)(1887,115){5}
wire [7:0] w58;    //: /sn:0 {0}(#:2132,448)(2012,448){1}
//: {2}(2008,448)(1629,448)(#:1629,217)(319,217){3}
//: {4}(317,215)(317,-520)(426,-520)(426,-569){5}
//: {6}(315,217)(226,217)(#:226,167){7}
//: {8}(2010,450)(2010,554)(2220,554){9}
wire [7:0] w65;    //: /sn:0 {0}(#:2132,401)(2123,401){1}
//: {2}(2119,401)(227,401)(#:227,344){3}
//: {4}(#:2121,403)(2121,507)(2220,507){5}
wire [7:0] w7;    //: /sn:0 {0}(#:1211,551)(1211,562)(1387,562)(1387,47)(1743,47){1}
//: {2}(1747,47)(1801,47){3}
//: {4}(1745,49)(1745,128)(1887,128){5}
wire w50;    //: /sn:0 {0}(-454,-238)(633,-238)(633,-196){1}
wire w59;    //: /sn:0 {0}(-548,-247)(-548,-228)(-483,-228){1}
wire w39;    //: /sn:0 {0}(232,-468)(232,-452)(118,-452)(118,-3){1}
//: {2}(120,-1)(203,-1){3}
//: {4}(118,1)(118,153)(135,153){5}
wire [7:0] w62;    //: /sn:0 {0}(2441,71)(2194,71)(2194,425)(#:2161,425){1}
wire [2:0] w4;    //: /sn:0 {0}(#:-615,-247)(-615,-174){1}
//: {2}(-613,-172)(620,-172){3}
//: {4}(-615,-170)(-615,-118)(-257,-118){5}
wire [7:0] w25;    //: /sn:0 {0}(#:1801,61)(1721,61){1}
//: {2}(1717,61)(1408,61)(1408,758)(1210,758)(#:1210,748){3}
//: {4}(1719,63)(1719,142)(1887,142){5}
wire [7:0] w56;    //: /sn:0 {0}(#:2132,435)(2045,435){1}
//: {2}(2041,435)(1517,435)(#:1517,803)(446,803)(#:446,748){3}
//: {4}(#:2043,437)(2043,541)(2220,541){5}
wire [7:0] w22;    //: /sn:0 {0}(#:226,12)(#:226,146){1}
wire w36;    //: /sn:0 {0}(954,540)(776,540)(776,-182)(649,-182){1}
wire [7:0] w0;    //: /sn:0 {0}(#:2132,421)(2076,421){1}
//: {2}(2072,421)(1554,421)(1554,608)(446,608)(#:446,551){3}
//: {4}(#:2074,423)(2074,527)(2220,527){5}
wire [7:0] w3;    //: /sn:0 {0}(445,146)(#:445,19){1}
wire w20;    //: /sn:0 {0}(909,152)(909,156)(953,156){1}
wire [7:0] Flag_shadow_output;    //: /sn:0 {0}(#:1125,-542)(1125,-487)(1326,-487)(1326,178){1}
//: {2}(1328,180)(1435,180)(1435,67)(1704,67){3}
//: {4}(1708,67)(1801,67){5}
//: {6}(1706,69)(1706,148)(1887,148){7}
//: {8}(1324,180)(1210,180)(#:1210,167){9}
wire w30;    //: /sn:0 {0}(897,-569)(897,-467)(385,-467)(385,4){1}
//: {2}(387,6)(422,6){3}
//: {4}(385,8)(385,94){5}
wire [7:0] w71;    //: /sn:0 {0}(#:990,167)(990,188)(1051,188){1}
//: {2}(1055,188)(1448,188)(1448,74)(1688,74){3}
//: {4}(1692,74)(1801,74){5}
//: {6}(1690,76)(1690,155)(1887,155){7}
//: {8}(1053,186)(1053,-517)(446,-517)(446,-569){9}
wire w42;    //: /sn:0 {0}(1173,737)(1157,737)(1157,699)(715,699)(715,-162)(649,-162){1}
wire [7:0] w37;    //: /sn:0 {0}(#:1801,27)(1794,27){1}
//: {2}(1790,27)(1376,27)(1376,365)(991,365)(#:991,344){3}
//: {4}(#:1792,29)(1792,108)(1887,108){5}
wire [7:0] w73;    //: /sn:0 {0}(#:1916,132)(2616,132)(2616,245)(2631,245){1}
wire w19;    //: /sn:0 {0}(-228,-108)(-176,-108)(-176,698)(396,698)(396,737)(409,737){1}
wire w12;    //: /sn:0 {0}(649,-155)(1115,-155)(1115,96)(1144,96)(1144,120){1}
wire [7:0] w18;    //: /sn:0 {0}(#:2132,415)(2090,415){1}
//: {2}(2086,415)(1565,415)(#:1565,617)(227,617)(#:227,551){3}
//: {4}(#:2088,417)(2088,521)(2220,521){5}
wire w23;    //: /sn:0 {0}(380,94)(380,86)(361,86)(361,-101)(-228,-101){1}
wire [7:0] w10;    //: /sn:0 {0}(#:1801,54)(1732,54){1}
//: {2}(1728,54)(1420,54)(1420,770)(991,770)(#:991,748){3}
//: {4}(1730,56)(1730,135)(1887,135){5}
wire [7:0] w84;    //: /sn:0 {0}(#:2249,531)(2616,531)(2616,265)(2631,265){1}
wire w24;    //: /sn:0 {0}(382,115)(382,156)(408,156){1}
wire w21;    //: /sn:0 {0}(156,156)(189,156){1}
wire w31;    //: /sn:0 {0}(954,333)(833,333)(833,-195)(649,-195){1}
wire [7:0] w1;    //: /sn:0 {0}(#:2132,428)(2059,428){1}
//: {2}(2055,428)(1530,428)(#:1530,813)(227,813)(#:227,748){3}
//: {4}(#:2057,430)(2057,534)(2220,534){5}
wire w32;    //: /sn:0 {0}(1771,-194)(1771,-183)(2647,-183)(2647,232){1}
wire w46;    //: /sn:0 {0}(1187,6)(1151,6){1}
//: {2}(1147,6)(1132,6)(1132,-466)(917,-466)(917,-569){3}
//: {4}(1149,8)(1149,120){5}
wire [7:0] w8;    //: /sn:0 {0}(1210,146)(#:1210,19){1}
wire w44;    //: /sn:0 {0}(252,-468)(252,-431)(912,-431)(912,-2){1}
//: {2}(914,0)(967,0){3}
//: {4}(912,2)(912,131){5}
wire w17;    //: /sn:0 {0}(649,-148)(879,-148)(879,102)(907,102)(907,131){1}
wire w27;    //: /sn:0 {0}(1684,-146)(1684,-119)(2457,-119)(2457,38){1}
wire [7:0] w28;    //: /sn:0 {0}(#:990,13)(#:990,146){1}
wire w35;    //: /sn:0 {0}(1174,540)(1154,540)(1154,499)(753,499)(753,-175)(649,-175){1}
wire w33;    //: /sn:0 {0}(1173,333)(1154,333)(1154,289)(798,289)(798,-188)(649,-188){1}
wire [7:0] w49;    //: /sn:0 {0}(2441,51)(#:1830,51){1}
wire w14;    //: /sn:0 {0}(-228,-134)(-6,-134)(-6,296)(399,296)(399,333)(409,333){1}
wire w45;    //: /sn:0 {0}(-33,-300)(335,-300){1}
//: {2}(339,-300)(532,-300){3}
//: {4}(536,-300)(1086,-300){5}
//: {6}(1090,-300)(1295,-300)(1295,149){7}
//: {8}(1293,151)(1249,151){9}
//: {10}(1295,153)(1295,326){11}
//: {12}(1293,328)(1249,328){13}
//: {14}(1295,330)(1295,533){15}
//: {16}(1293,535)(1250,535){17}
//: {18}(1295,537)(1295,732)(1249,732){19}
//: {20}(1088,-298)(1088,149){21}
//: {22}(1086,151)(1029,151){23}
//: {24}(1088,153)(1088,326){25}
//: {26}(1086,328)(1030,328){27}
//: {28}(1088,330)(1088,533){29}
//: {30}(1086,535)(1030,535){31}
//: {32}(1088,537)(1088,732)(1030,732){33}
//: {34}(534,-298)(534,149){35}
//: {36}(532,151)(484,151){37}
//: {38}(534,153)(534,326){39}
//: {40}(532,328)(485,328){41}
//: {42}(534,330)(534,533){43}
//: {44}(532,535)(485,535){45}
//: {46}(534,537)(534,732)(485,732){47}
//: {48}(337,-298)(337,149){49}
//: {50}(335,151)(265,151){51}
//: {52}(337,153)(337,326){53}
//: {54}(335,328)(266,328){55}
//: {56}(337,330)(337,533){57}
//: {58}(335,535)(266,535){59}
//: {60}(337,537)(337,732)(266,732){61}
wire w2;    //: /sn:0 {0}(-228,-141)(28,-141)(28,333)(190,333){1}
wire w41;    //: /sn:0 {0}(190,540)(-77,540)(-77,-128)(-228,-128){1}
wire w11;    //: /sn:0 {0}(1173,156)(1146,156)(1146,141){1}
wire w47;    //: /sn:0 {0}(190,737)(-161,737)(-161,-114)(-228,-114){1}
wire [7:0] w15;    //: /sn:0 {0}(#:1105,-542)(1105,-447)(507,-447)(507,205){1}
//: {2}(509,207)(1640,207)(1640,441)(2025,441){3}
//: {4}(2029,441)(2132,441){5}
//: {6}(2027,443)(2027,547)(2220,547){7}
//: {8}(505,207)(445,207)(#:445,167){9}
wire [2:0] w83;    //: /sn:0 {0}(#:2236,508)(2236,-80)(1905,-80){1}
//: {2}(1901,-80)(1740,-80)(#:1740,-194){3}
//: {4}(1903,-78)(1903,109){5}
wire [2:0] w5;    //: /sn:0 {0}(#:1817,28)(1817,-22){1}
//: {2}(#:1819,-24)(2148,-24)(2148,402){3}
//: {4}(1815,-24)(1656,-24)(#:1656,-146){5}
wire w38;    //: /sn:0 {0}(409,540)(389,540)(389,494)(-110,494)(-110,-121)(-228,-121){1}
wire w43;    //: /sn:0 {0}(954,737)(735,737)(735,-168)(649,-168){1}
wire w9;    //: /sn:0 {0}(-454,-218)(-244,-218)(-244,-142){1}
wire w26;    //: /sn:0 {0}(-228,-94)(105,-94)(105,158)(135,158){1}
//: enddecls

  //: IN g116 (Accumulator_input) @(216,-403) /sn:0 /R:3 /w:[ 0 ]
  //: joint g4 (w80) @(613, 545) /w:[ -1 18 24 17 ]
  //: joint g8 (w80) @(1278, 742) /w:[ -1 34 44 33 ]
  //: joint g17 (w80) @(300, 338) /w:[ -1 1 2 4 ]
  _GGREG8 #(10, 10, 20) C0 (.Q(w6), .D(Register_input), .EN(w80), .CLR(w45), .CK(w33));   //: @(1210,333) /w:[ 0 25 41 13 0 ]
  //: joint g74 (w7) @(1745, 47) /w:[ 2 -1 1 4 ]
  //: joint g30 (w45) @(1295, 151) /w:[ -1 7 8 10 ]
  //: joint g92 (w46) @(1149, 6) /w:[ 1 -1 2 4 ]
  //: joint g77 (w25) @(1719, 61) /w:[ 1 -1 2 4 ]
  //: frame g1 @(923,110) /sn:0 /wi:391 /ht:679 /tx:"Shadow registers"
  //: joint g111 (Use_shadow_reg) @(656, -558) /w:[ 2 4 -1 1 ]
  _GGREG8 #(10, 10, 20) A (.Q(w58), .D(w22), .EN(w80), .CLR(w45), .CK(w21));   //: @(226,156) /w:[ 7 1 0 51 1 ]
  //: OUT g51 (Register_output2) @(2814,254) /sn:0 /w:[ 1 ]
  //: joint g70 (w16) @(1761, 41) /w:[ 2 -1 1 4 ]
  //: joint g103 (w15) @(2027, 441) /w:[ 4 -1 3 6 ]
  //: joint g10 (w80) @(1278, 338) /w:[ -1 38 40 37 ]
  //: joint g25 (w45) @(1088, 535) /w:[ -1 29 30 32 ]
  //: joint g65 (Flag_shadow_output) @(1326, 180) /w:[ 2 1 8 -1 ]
  //: joint g64 (w5) @(1817, -24) /w:[ 2 -1 4 1 ]
  //: IN g72 (Register_output_choose2) @(1630,-198) /sn:0 /w:[ 0 ]
  //: joint g49 (Register_input) @(991, 518) /w:[ 40 -1 39 42 ]
  //: joint g6 (w80) @(613, 861) /w:[ 30 29 -1 60 ]
  //: joint g35 (Register_input) @(-340, -52) /w:[ 2 -1 1 16 ]
  //: joint g7 (w80) @(1066, 861) /w:[ 32 46 31 -1 ]
  assign w4 = Register_input_choose[2:0]; //: TAP g56 @(-615,-253) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g58 (w4) @(-615, -172) /w:[ 2 1 -1 4 ]
  //: joint g98 (w13) @(2104, 408) /w:[ 1 -1 2 4 ]
  //: joint g85 (Flag_shadow_output) @(1706, 67) /w:[ 4 -1 3 6 ]
  //: joint g67 (w83) @(1903, -80) /w:[ 1 -1 2 4 ]
  //: joint g33 (w45) @(534, -300) /w:[ 4 -1 3 34 ]
  //: joint g54 (w45) @(337, -300) /w:[ 2 -1 1 48 ]
  //: joint g81 (Flag_input) @(760, -383) /w:[ 1 2 4 -1 ]
  //: joint g40 (Register_input) @(446, 311) /w:[ 22 -1 21 28 ]
  _GGDECODER8 #(6, 6) g52 (.I(w4), .E(w9), .Z0(w2), .Z1(w14), .Z2(w41), .Z3(w38), .Z4(w47), .Z5(w19), .Z6(w23), .Z7(w26));   //: @(-244,-118) /sn:0 /R:1 /w:[ 5 1 0 0 1 1 1 0 1 0 ] /ss:1 /do:1
  assign w32 = Register_output_choose2[3]; //: TAP g108 @(1771,-200) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g12 (w80) @(1066, 545) /w:[ -1 50 56 49 ]
  _GGMUX2x8 #(8, 8) g106 (.I0(w84), .I1(w73), .S(w32), .Z(Register_output2));   //: @(2647,255) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:1 /do:0
  _GGREG8 #(10, 10, 20) H0 (.Q(w10), .D(Register_input), .EN(w80), .CLR(w45), .CK(w43));   //: @(991,737) /w:[ 3 57 59 33 0 ]
  assign w83 = Register_output_choose2[2:0]; //: TAP g96 @(1740,-200) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  //: joint g117 (Accumulator_input) @(216, -330) /w:[ 2 1 -1 4 ]
  //: joint g114 (Register_input) @(1000, -52) /w:[ 8 -1 7 10 ]
  _GGREG8 #(10, 10, 20) C (.Q(w13), .D(Register_input), .EN(w80), .CLR(w45), .CK(w14));   //: @(446,333) /w:[ 3 29 23 41 1 ]
  _GGREG8 #(10, 10, 20) D (.Q(w18), .D(Register_input), .EN(w80), .CLR(w45), .CK(w41));   //: @(227,540) /w:[ 3 47 7 59 0 ]
  //: joint g19 (w45) @(534, 535) /w:[ -1 43 44 46 ]
  //: OUT g78 (Flag_output) @(1115,-651) /sn:0 /R:1 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) L0 (.Q(w25), .D(Register_input), .EN(w80), .CLR(w45), .CK(w42));   //: @(1210,737) /w:[ 3 55 45 19 0 ]
  //: joint g113 (w44) @(912, 0) /w:[ 2 1 -1 4 ]
  _GGMUX2x8 #(8, 8) g105 (.I0(w62), .I1(w49), .S(w27), .Z(Register_output1));   //: @(2457,61) /sn:0 /R:1 /w:[ 0 0 1 0 ] /ss:1 /do:0
  //: joint g100 (w0) @(2074, 421) /w:[ 1 -1 2 4 ]
  assign w5 = Register_output_choose1[2:0]; //: TAP g93 @(1656,-152) /sn:0 /R:1 /w:[ 5 1 2 ] /ss:1
  _GGMUX8x8 #(20, 20) g63 (.I0(w65), .I1(w13), .I2(w18), .I3(w0), .I4(w1), .I5(w56), .I6(w15), .I7(w58), .S(w83), .Z(w84));   //: @(2236,531) /sn:0 /R:1 /w:[ 5 5 5 5 5 5 7 9 0 0 ] /ss:1 /do:1
  _GGMUX2x8 #(8, 8) g38 (.I0(Register_input), .I1(Accumulator_input), .S(w39), .Z(w22));   //: @(226,-1) /sn:0 /w:[ 15 5 3 0 ] /ss:0 /do:1
  //: joint g101 (w1) @(2057, 428) /w:[ 1 -1 2 4 ]
  //: frame g0 @(150,111) /sn:0 /wi:399 /ht:676 /tx:"Main registers"
  //: joint g43 (Register_input) @(-340, 518) /w:[ 34 33 -1 48 ]
  //: joint g48 (Register_input) @(446, 518) /w:[ 38 -1 37 44 ]
  _GGMUX2x8 #(8, 8) g37 (.I0(Register_input), .I1(Flag_input), .S(w30), .Z(w3));   //: @(445,6) /sn:0 /w:[ 13 5 3 1 ] /ss:0 /do:1
  //: joint g122 (w58) @(317, 217) /w:[ 3 4 6 -1 ]
  //: comment g120 @(1436,4) /sn:0
  //: /line:"Shadow regs"
  //: /end
  //: joint g95 (w71) @(1690, 74) /w:[ 4 -1 3 6 ]
  //: IN g80 (Flag_input) @(760,-401) /sn:0 /R:3 /w:[ 3 ]
  _GGREG8 #(10, 10, 20) B0 (.Q(w37), .D(Register_input), .EN(w80), .CLR(w45), .CK(w31));   //: @(991,333) /w:[ 3 27 55 27 0 ]
  //: joint g76 (w10) @(1730, 54) /w:[ 1 -1 2 4 ]
  _GGREG8 #(10, 10, 20) A0 (.Q(w71), .D(w28), .EN(w80), .CLR(w45), .CK(w20));   //: @(990,156) /w:[ 0 1 53 23 1 ]
  //: joint g44 (Register_input) @(227, 716) /w:[ 50 -1 49 60 ]
  //: VDD g75 (w40) @(-459,-295) /sn:0 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) B (.Q(w65), .D(Register_input), .EN(w80), .CLR(w45), .CK(w2));   //: @(227,333) /w:[ 3 31 3 55 1 ]
  //: joint g3 (w80) @(613, 742) /w:[ -1 16 26 15 ]
  //: joint g16 (w80) @(300, 742) /w:[ -1 9 10 12 ]
  //: joint g47 (Register_input) @(227, 518) /w:[ 36 -1 35 46 ]
  _GGMUX2x8 #(8, 8) g109 (.I0(w15), .I1(Flag_shadow_output), .S(Use_shadow_reg), .Z(Flag_output));   //: @(1115,-558) /sn:0 /R:2 /w:[ 0 0 3 1 ] /ss:1 /do:1
  //: joint g26 (w45) @(1088, 328) /w:[ -1 25 26 28 ]
  _GGOR2 #(6) g90 (.I0(w39), .I1(w26), .Z(w21));   //: @(146,156) /sn:0 /w:[ 5 1 0 ]
  //: GROUND g2 (w80) @(613,931) /sn:0 /w:[ 61 ]
  _GGREG8 #(10, 10, 20) F (.Q(w15), .D(w3), .EN(w80), .CLR(w45), .CK(w24));   //: @(445,156) /w:[ 9 0 21 37 1 ]
  //: joint g23 (w45) @(337, 535) /w:[ -1 57 58 60 ]
  _GGOR2 #(6) g91 (.I0(w46), .I1(w12), .Z(w11));   //: @(1146,131) /sn:0 /R:3 /w:[ 5 1 1 ]
  //: joint g104 (w58) @(2010, 448) /w:[ 1 -1 2 8 ]
  //: IN g86 (Flag_input_choose) @(907,-627) /sn:0 /R:3 /w:[ 1 ]
  //: joint g24 (w45) @(337, 328) /w:[ -1 53 54 56 ]
  //: joint g39 (Register_input) @(227, 311) /w:[ 20 -1 19 30 ]
  //: comment g121 @(1723,378) /sn:0
  //: /line:"Normal regs"
  //: /end
  //: joint g29 (w45) @(1295, 328) /w:[ -1 11 12 14 ]
  _GGMUX8x8 #(20, 20) g60 (.I0(w37), .I1(w6), .I2(w16), .I3(w7), .I4(w10), .I5(w25), .I6(Flag_shadow_output), .I7(w71), .S(w5), .Z(w49));   //: @(1817,51) /sn:0 /R:1 /w:[ 0 3 3 3 0 0 5 5 0 1 ] /ss:1 /do:1
  _GGDECODER2 #(6, 6) g110 (.I(Accumulator_input_choose), .E(Use_shadow_reg), .Z0(w39), .Z1(w44));   //: @(242,-484) /sn:0 /w:[ 1 0 0 0 ] /ss:1 /do:0
  _GGMUX2x8 #(8, 8) g82 (.I0(Register_input), .I1(Flag_input), .S(w46), .Z(w8));   //: @(1210,6) /sn:0 /w:[ 9 0 0 1 ] /ss:0 /do:1
  //: IN g18 (Register_reset) @(-66,-300) /sn:0 /w:[ 1 ]
  _GGMUX2x8 #(8, 8) g119 (.I0(w58), .I1(w71), .S(Use_shadow_reg), .Z(Accumulator_output));   //: @(436,-585) /sn:0 /R:2 /w:[ 5 9 11 0 ] /ss:0 /do:1
  _GGOR2 #(6) g94 (.I0(w30), .I1(w23), .Z(w24));   //: @(382,105) /sn:0 /R:3 /w:[ 5 0 0 ]
  assign w27 = Register_output_choose1[3]; //: TAP g107 @(1684,-152) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  _GGREG8 #(10, 10, 20) E0 (.Q(w7), .D(Register_input), .EN(w80), .CLR(w45), .CK(w35));   //: @(1211,540) /w:[ 0 41 43 17 0 ]
  _GGREG8 #(10, 10, 20) D0 (.Q(w16), .D(Register_input), .EN(w80), .CLR(w45), .CK(w36));   //: @(991,540) /w:[ 0 43 57 31 0 ]
  //: OUT g50 (Register_output1) @(2814,61) /sn:0 /w:[ 1 ]
  //: joint g9 (w80) @(1278, 545) /w:[ -1 36 42 35 ]
  //: IN g73 (Register_input_choose) @(-673,-251) /sn:0 /w:[ 0 ]
  //: joint g68 (w37) @(1792, 27) /w:[ 1 -1 2 4 ]
  //: joint g102 (w56) @(2043, 435) /w:[ 1 -1 2 4 ]
  //: IN g71 (Register_output_choose1) @(1576,-150) /sn:0 /w:[ 0 ]
  //: joint g22 (w45) @(337, 151) /w:[ -1 49 50 52 ]
  _GGNBUF #(2) g31 (.I(Register_reset), .Z(w45));   //: @(-43,-300) /sn:0 /w:[ 0 0 ]
  //: joint g59 (w30) @(385, 6) /w:[ 2 1 -1 4 ]
  _GGDECODER2 #(6, 6) g87 (.I(Flag_input_choose), .E(Use_shadow_reg), .Z0(w30), .Z1(w46));   //: @(907,-585) /sn:0 /w:[ 0 7 0 3 ] /ss:0 /do:0
  _GGMUX2x8 #(8, 8) g83 (.I0(Register_input), .I1(Accumulator_input), .S(w44), .Z(w28));   //: @(990,0) /sn:0 /w:[ 11 3 3 0 ] /ss:0 /do:1
  //: joint g99 (w18) @(2088, 415) /w:[ 1 -1 2 4 ]
  //: joint g45 (Register_input) @(446, 716) /w:[ 52 -1 51 58 ]
  //: joint g41 (Register_input) @(991, 311) /w:[ 24 -1 23 26 ]
  _GGOR2 #(6) g36 (.I0(w44), .I1(w17), .Z(w20));   //: @(909,142) /sn:0 /R:3 /w:[ 5 1 0 ]
  //: joint g42 (Register_input) @(-340, 311) /w:[ 18 17 -1 32 ]
  //: joint g69 (w6) @(1776, 34) /w:[ 2 -1 1 4 ]
  //: joint g66 (w15) @(507, 207) /w:[ 2 1 8 -1 ]
  //: joint g28 (w45) @(1295, 535) /w:[ -1 15 16 18 ]
  //: IN g34 (Register_input) @(-388,-52) /sn:0 /w:[ 0 ]
  //: joint g46 (Register_input) @(991, 716) /w:[ 54 -1 53 56 ]
  assign w59 = Register_input_choose[3]; //: TAP g57 @(-548,-253) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: OUT g118 (Accumulator_output) @(436,-661) /sn:0 /R:1 /w:[ 1 ]
  //: joint g84 (Register_input) @(455, -52) /w:[ 6 -1 5 12 ]
  //: joint g5 (w80) @(613, 338) /w:[ -1 20 22 19 ]
  //: joint g11 (w80) @(1066, 338) /w:[ -1 52 54 51 ]
  //: joint g14 (w80) @(613, 854) /w:[ -1 14 13 28 ]
  //: joint g112 (w39) @(118, -1) /w:[ 2 1 -1 4 ]
  _GGREG8 #(10, 10, 20) H (.Q(w1), .D(Register_input), .EN(w80), .CLR(w45), .CK(w47));   //: @(227,737) /w:[ 3 61 11 61 0 ]
  //: joint g123 (w71) @(1053, 188) /w:[ 2 8 1 -1 ]
  //: joint g21 (w45) @(534, 151) /w:[ -1 35 36 38 ]
  _GGMUX8x8 #(20, 20) g61 (.I0(w65), .I1(w13), .I2(w18), .I3(w0), .I4(w1), .I5(w56), .I6(w15), .I7(w58), .S(w5), .Z(w62));   //: @(2148,425) /sn:0 /R:1 /w:[ 0 0 0 0 0 0 5 0 3 1 ] /ss:1 /do:1
  //: joint g115 (Register_input) @(236, -52) /w:[ 4 -1 3 14 ]
  //: joint g79 (Use_shadow_reg) @(656, -585) /w:[ 6 8 10 5 ]
  //: joint g20 (w45) @(534, 328) /w:[ -1 39 40 42 ]
  //: joint g32 (w45) @(1088, -300) /w:[ 6 -1 5 20 ]
  //: joint g97 (w65) @(2121, 401) /w:[ 1 -1 2 4 ]
  //: IN g89 (Use_shadow_reg) @(656,-624) /sn:0 /R:3 /w:[ 9 ]
  //: joint g15 (w80) @(300, 545) /w:[ -1 5 6 8 ]
  _GGREG8 #(10, 10, 20) E (.Q(w0), .D(Register_input), .EN(w80), .CLR(w45), .CK(w38));   //: @(446,540) /w:[ 3 45 25 45 0 ]
  //: joint g27 (w45) @(1088, 151) /w:[ -1 21 22 24 ]
  _GGREG8 #(10, 10, 20) F0 (.Q(Flag_shadow_output), .D(w8), .EN(w80), .CLR(w45), .CK(w11));   //: @(1210,156) /w:[ 9 0 39 9 0 ]
  _GGMUX8x8 #(20, 20) g62 (.I0(w37), .I1(w6), .I2(w16), .I3(w7), .I4(w10), .I5(w25), .I6(Flag_shadow_output), .I7(w71), .S(w83), .Z(w73));   //: @(1903,132) /sn:0 /R:1 /w:[ 5 5 5 5 5 5 7 7 5 0 ] /ss:1 /do:1
  //: IN g88 (Accumulator_input_choose) @(197,-651) /sn:0 /R:3 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) L (.Q(w56), .D(Register_input), .EN(w80), .CLR(w45), .CK(w19));   //: @(446,737) /w:[ 3 59 27 47 1 ]
  _GGDECODER2 #(6, 6) g55 (.I(w59), .E(w40), .Z0(w9), .Z1(w50));   //: @(-470,-228) /sn:0 /R:1 /w:[ 1 1 0 0 ] /ss:1 /do:0
  //: joint g13 (w80) @(1066, 742) /w:[ -1 48 58 47 ]
  _GGDECODER8 #(6, 6) g53 (.I(w4), .E(w50), .Z0(w31), .Z1(w33), .Z2(w36), .Z3(w35), .Z4(w43), .Z5(w42), .Z6(w12), .Z7(w17));   //: @(633,-172) /sn:0 /R:1 /w:[ 3 1 1 1 1 1 1 1 0 0 ] /ss:1 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin instruction_IX
module instruction_IX(CB, Instruction_input);
//: interface  /sz:(303, 522) /bd:[ Li0>Instruction_input[7:0](208/522) Bo0<CB(20/303) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
output CB;    //: /sn:0 {0}(-106,580)(636,580)(636,306){1}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire w139;    //: /sn:0 {0}(924,306)(924,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire w128;    //: /sn:0 {0}(963,306)(963,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w86;    //: /sn:0 {0}(633,306)(633,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,321){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w140;    //: /sn:0 {0}(921,306)(921,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w147;    //: /sn:0 {0}(1049,306)(1049,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w260;    //: /sn:0 {0}(1571,306)(1571,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w44;    //: /sn:0 {0}(464,306)(464,321){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w135;    //: /sn:0 {0}(938,306)(938,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w11;    //: /sn:0 {0}(254,218)(898,218)(898,290)(913,290){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,321){1}
wire w129;    //: /sn:0 {0}(959,306)(959,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w286;    //: /sn:0 {0}(1624,306)(1624,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w158;    //: /sn:0 {0}(1011,306)(1011,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w142;    //: /sn:0 {0}(914,306)(914,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w148;    //: /sn:0 {0}(1046,306)(1046,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w154;    //: /sn:0 {0}(1025,306)(1025,321){1}
wire w156;    //: /sn:0 {0}(1018,306)(1018,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w130;    //: /sn:0 {0}(956,306)(956,321){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w131;    //: /sn:0 {0}(952,306)(952,321){1}
wire w268;    //: /sn:0 {0}(1543,306)(1543,321){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w304;    //: /sn:0 {0}(1703,306)(1703,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w52;    //: /sn:0 {0}(436,306)(436,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w150;    //: /sn:0 {0}(1039,306)(1039,321){1}
wire w33;    //: /sn:0 {0}(343,306)(343,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w69;    //: /sn:0 {0}(540,306)(540,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w146;    //: /sn:0 {0}(1053,306)(1053,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w151;    //: /sn:0 {0}(1035,306)(1035,321){1}
wire w161;    //: /sn:0 {0}(1000,306)(1000,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w137;    //: /sn:0 {0}(931,306)(931,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w157;    //: /sn:0 {0}(1014,306)(1014,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w132;    //: /sn:0 {0}(949,306)(949,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w152;    //: /sn:0 {0}(1032,306)(1032,321){1}
wire w138;    //: /sn:0 {0}(928,306)(928,321){1}
wire w269;    //: /sn:0 {0}(1539,306)(1539,321){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w136;    //: /sn:0 {0}(935,306)(935,321){1}
wire w134;    //: /sn:0 {0}(942,306)(942,321){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w153;    //: /sn:0 {0}(1028,306)(1028,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w155;    //: /sn:0 {0}(1021,306)(1021,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w26;    //: /sn:0 {0}(368,306)(368,321){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w143;    //: /sn:0 {0}(910,306)(910,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w278;    //: /sn:0 {0}(1652,306)(1652,321){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w159;    //: /sn:0 {0}(1007,306)(1007,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w141;    //: /sn:0 {0}(917,306)(917,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w10;    //: /sn:0 {0}(254,214)(988,214)(988,290)(1003,290){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(935,156){13}
//: {14}(#:939,156)(1025,156){15}
//: {16}(#:1029,156)(1118,156){17}
//: {18}(#:1122,156)(1208,156){19}
//: {20}(#:1212,156)(1297,156){21}
//: {22}(#:1301,156)(1391,156){23}
//: {24}(#:1395,156)(1481,156){25}
//: {26}(#:1485,156)(1564,156){27}
//: {28}(#:1568,156)(1645,156){29}
//: {30}(#:1649,156)(1726,156)(1726,277){31}
//: {32}(1647,158)(1647,277){33}
//: {34}(1566,158)(1566,277){35}
//: {36}(1483,158)(1483,277){37}
//: {38}(1393,158)(1393,277){39}
//: {40}(1299,158)(1299,277){41}
//: {42}(1210,158)(1210,277){43}
//: {44}(1120,158)(1120,277){45}
//: {46}(1027,158)(1027,277){47}
//: {48}(937,158)(937,277){49}
//: {50}(842,158)(842,277){51}
//: {52}(744,158)(744,277){53}
//: {54}(649,158)(649,277){55}
//: {56}(560,158)(560,277){57}
//: {58}(459,158)(459,277){59}
//: {60}(363,158)(363,277){61}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w290;    //: /sn:0 {0}(1752,306)(1752,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w80;    //: /sn:0 {0}(654,306)(654,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire w277;    //: /sn:0 {0}(1655,306)(1655,321){1}
wire w149;    //: /sn:0 {0}(1042,306)(1042,321){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w160;    //: /sn:0 {0}(1004,306)(1004,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire w133;    //: /sn:0 {0}(945,306)(945,321){1}
wire w77;    //: /sn:0 {0}(664,306)(664,321){1}
wire w51;    //: /sn:0 {0}(439,306)(439,321){1}
//: enddecls

  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 53 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(w26), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(w33), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 61 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 37 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 50 ]
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(w269));   //: @(1566,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w1) @(1210, 156) /w:[ 20 -1 19 42 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 56 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 54 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g29 (w1) @(1120, 156) /w:[ 18 -1 17 44 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 52 ]
  _GGDECODER16 #(6, 6) g10 (.I(w1), .E(w11), .Z0(w128), .Z1(w129), .Z2(w130), .Z3(w131), .Z4(w132), .Z5(w133), .Z6(w134), .Z7(w135), .Z8(w136), .Z9(w137), .Z10(w138), .Z11(w139), .Z12(w140), .Z13(w141), .Z14(w142), .Z15(w143));   //: @(937,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(w69), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 57 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 30 -1 29 32 ]
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 51 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(w77), .Z4(w78), .Z5(w79), .Z6(w80), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(CB), .Z12(w86), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 55 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w1) @(1299, 156) /w:[ 22 -1 21 40 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 58 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: joint g33 (w1) @(1483, 156) /w:[ 26 -1 25 36 ]
  //: OUT g40 (CB) @(-103,580) /sn:0 /R:2 /w:[ 0 ]
  _GGDECODER16 #(6, 6) g12 (.I(w1), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g34 (w1) @(1566, 156) /w:[ 28 -1 27 34 ]
  //: joint g28 (w1) @(1027, 156) /w:[ 16 -1 15 46 ]
  _GGDECODER16 #(6, 6) g14 (.I(w1), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g11 (.I(w1), .E(w10), .Z0(w146), .Z1(w147), .Z2(w148), .Z3(w149), .Z4(w150), .Z5(w151), .Z6(w152), .Z7(w153), .Z8(w154), .Z9(w155), .Z10(w156), .Z11(w157), .Z12(w158), .Z13(w159), .Z14(w160), .Z15(w161));   //: @(1027,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(w44), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(w51), .Z14(w52), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 59 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 60 ]
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(w290), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 31 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g32 (w1) @(1393, 156) /w:[ 24 -1 23 38 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w1), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: joint g27 (w1) @(937, 156) /w:[ 14 -1 13 48 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w1), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 43 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin instruction_BITS
module instruction_BITS(Instruction_input);
//: interface  /sz:(317, 550) /bd:[ Li0>Instruction_input[7:0](220/550) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire w139;    //: /sn:0 {0}(924,306)(924,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire w128;    //: /sn:0 {0}(963,306)(963,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w86;    //: /sn:0 {0}(633,306)(633,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,321){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w140;    //: /sn:0 {0}(921,306)(921,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w147;    //: /sn:0 {0}(1049,306)(1049,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w260;    //: /sn:0 {0}(1571,306)(1571,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w44;    //: /sn:0 {0}(464,306)(464,321){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w135;    //: /sn:0 {0}(938,306)(938,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w11;    //: /sn:0 {0}(254,218)(898,218)(898,290)(913,290){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,321){1}
wire w129;    //: /sn:0 {0}(959,306)(959,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w286;    //: /sn:0 {0}(1624,306)(1624,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w158;    //: /sn:0 {0}(1011,306)(1011,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w142;    //: /sn:0 {0}(914,306)(914,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w148;    //: /sn:0 {0}(1046,306)(1046,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w154;    //: /sn:0 {0}(1025,306)(1025,321){1}
wire w156;    //: /sn:0 {0}(1018,306)(1018,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w130;    //: /sn:0 {0}(956,306)(956,321){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w131;    //: /sn:0 {0}(952,306)(952,321){1}
wire w268;    //: /sn:0 {0}(1543,306)(1543,321){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w304;    //: /sn:0 {0}(1703,306)(1703,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w52;    //: /sn:0 {0}(436,306)(436,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w150;    //: /sn:0 {0}(1039,306)(1039,321){1}
wire w33;    //: /sn:0 {0}(343,306)(343,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w69;    //: /sn:0 {0}(540,306)(540,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w146;    //: /sn:0 {0}(1053,306)(1053,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w85;    //: /sn:0 {0}(636,306)(636,321){1}
wire w151;    //: /sn:0 {0}(1035,306)(1035,321){1}
wire w161;    //: /sn:0 {0}(1000,306)(1000,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w137;    //: /sn:0 {0}(931,306)(931,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w157;    //: /sn:0 {0}(1014,306)(1014,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w132;    //: /sn:0 {0}(949,306)(949,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w152;    //: /sn:0 {0}(1032,306)(1032,321){1}
wire w138;    //: /sn:0 {0}(928,306)(928,321){1}
wire w269;    //: /sn:0 {0}(1539,306)(1539,321){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w136;    //: /sn:0 {0}(935,306)(935,321){1}
wire w134;    //: /sn:0 {0}(942,306)(942,321){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w153;    //: /sn:0 {0}(1028,306)(1028,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w155;    //: /sn:0 {0}(1021,306)(1021,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w26;    //: /sn:0 {0}(368,306)(368,321){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w143;    //: /sn:0 {0}(910,306)(910,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w278;    //: /sn:0 {0}(1652,306)(1652,321){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w159;    //: /sn:0 {0}(1007,306)(1007,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w141;    //: /sn:0 {0}(917,306)(917,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w10;    //: /sn:0 {0}(254,214)(988,214)(988,290)(1003,290){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(935,156){13}
//: {14}(#:939,156)(1025,156){15}
//: {16}(#:1029,156)(1118,156){17}
//: {18}(#:1122,156)(1208,156){19}
//: {20}(#:1212,156)(1297,156){21}
//: {22}(#:1301,156)(1391,156){23}
//: {24}(#:1395,156)(1481,156){25}
//: {26}(#:1485,156)(1564,156){27}
//: {28}(#:1568,156)(1645,156){29}
//: {30}(#:1649,156)(1726,156)(1726,277){31}
//: {32}(1647,158)(1647,277){33}
//: {34}(1566,158)(1566,277){35}
//: {36}(1483,158)(1483,277){37}
//: {38}(1393,158)(1393,277){39}
//: {40}(1299,158)(1299,277){41}
//: {42}(1210,158)(1210,277){43}
//: {44}(1120,158)(1120,277){45}
//: {46}(1027,158)(1027,277){47}
//: {48}(937,158)(937,277){49}
//: {50}(842,158)(842,277){51}
//: {52}(744,158)(744,277){53}
//: {54}(649,158)(649,277){55}
//: {56}(560,158)(560,277){57}
//: {58}(459,158)(459,277){59}
//: {60}(363,158)(363,277){61}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w290;    //: /sn:0 {0}(1752,306)(1752,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w80;    //: /sn:0 {0}(654,306)(654,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire w277;    //: /sn:0 {0}(1655,306)(1655,321){1}
wire w149;    //: /sn:0 {0}(1042,306)(1042,321){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w160;    //: /sn:0 {0}(1004,306)(1004,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire w133;    //: /sn:0 {0}(945,306)(945,321){1}
wire w77;    //: /sn:0 {0}(664,306)(664,321){1}
wire w51;    //: /sn:0 {0}(439,306)(439,321){1}
//: enddecls

  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 53 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(w26), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(w33), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 61 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 37 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 50 ]
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(w269));   //: @(1566,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w1) @(1210, 156) /w:[ 20 -1 19 42 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 56 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 54 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g29 (w1) @(1120, 156) /w:[ 18 -1 17 44 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 52 ]
  _GGDECODER16 #(6, 6) g10 (.I(w1), .E(w11), .Z0(w128), .Z1(w129), .Z2(w130), .Z3(w131), .Z4(w132), .Z5(w133), .Z6(w134), .Z7(w135), .Z8(w136), .Z9(w137), .Z10(w138), .Z11(w139), .Z12(w140), .Z13(w141), .Z14(w142), .Z15(w143));   //: @(937,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(w69), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 57 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 30 -1 29 32 ]
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 51 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(w77), .Z4(w78), .Z5(w79), .Z6(w80), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(w85), .Z12(w86), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 55 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w1) @(1299, 156) /w:[ 22 -1 21 40 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 58 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: joint g33 (w1) @(1483, 156) /w:[ 26 -1 25 36 ]
  _GGDECODER16 #(6, 6) g12 (.I(w1), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g34 (w1) @(1566, 156) /w:[ 28 -1 27 34 ]
  //: joint g28 (w1) @(1027, 156) /w:[ 16 -1 15 46 ]
  _GGDECODER16 #(6, 6) g14 (.I(w1), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g11 (.I(w1), .E(w10), .Z0(w146), .Z1(w147), .Z2(w148), .Z3(w149), .Z4(w150), .Z5(w151), .Z6(w152), .Z7(w153), .Z8(w154), .Z9(w155), .Z10(w156), .Z11(w157), .Z12(w158), .Z13(w159), .Z14(w160), .Z15(w161));   //: @(1027,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(w44), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(w51), .Z14(w52), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 59 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 60 ]
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(w290), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 31 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g32 (w1) @(1393, 156) /w:[ 24 -1 23 38 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w1), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: joint g27 (w1) @(937, 156) /w:[ 14 -1 13 48 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w1), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 43 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin instruction_IX_BITS
module instruction_IX_BITS(Instruction_input);
//: interface  /sz:(333, 562) /bd:[ Li0>Instruction_input[7:0](224/562) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire w139;    //: /sn:0 {0}(924,306)(924,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire w128;    //: /sn:0 {0}(963,306)(963,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w86;    //: /sn:0 {0}(633,306)(633,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,321){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w140;    //: /sn:0 {0}(921,306)(921,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w147;    //: /sn:0 {0}(1049,306)(1049,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w260;    //: /sn:0 {0}(1571,306)(1571,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w44;    //: /sn:0 {0}(464,306)(464,321){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w135;    //: /sn:0 {0}(938,306)(938,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w11;    //: /sn:0 {0}(254,218)(898,218)(898,290)(913,290){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,321){1}
wire w129;    //: /sn:0 {0}(959,306)(959,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w286;    //: /sn:0 {0}(1624,306)(1624,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w158;    //: /sn:0 {0}(1011,306)(1011,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w142;    //: /sn:0 {0}(914,306)(914,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w148;    //: /sn:0 {0}(1046,306)(1046,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w154;    //: /sn:0 {0}(1025,306)(1025,321){1}
wire w156;    //: /sn:0 {0}(1018,306)(1018,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w130;    //: /sn:0 {0}(956,306)(956,321){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w131;    //: /sn:0 {0}(952,306)(952,321){1}
wire w268;    //: /sn:0 {0}(1543,306)(1543,321){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w304;    //: /sn:0 {0}(1703,306)(1703,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w52;    //: /sn:0 {0}(436,306)(436,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w150;    //: /sn:0 {0}(1039,306)(1039,321){1}
wire w33;    //: /sn:0 {0}(343,306)(343,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w69;    //: /sn:0 {0}(540,306)(540,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w146;    //: /sn:0 {0}(1053,306)(1053,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w85;    //: /sn:0 {0}(636,306)(636,321){1}
wire w151;    //: /sn:0 {0}(1035,306)(1035,321){1}
wire w161;    //: /sn:0 {0}(1000,306)(1000,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w137;    //: /sn:0 {0}(931,306)(931,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w157;    //: /sn:0 {0}(1014,306)(1014,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w132;    //: /sn:0 {0}(949,306)(949,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w152;    //: /sn:0 {0}(1032,306)(1032,321){1}
wire w138;    //: /sn:0 {0}(928,306)(928,321){1}
wire w269;    //: /sn:0 {0}(1539,306)(1539,321){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w136;    //: /sn:0 {0}(935,306)(935,321){1}
wire w134;    //: /sn:0 {0}(942,306)(942,321){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w153;    //: /sn:0 {0}(1028,306)(1028,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w155;    //: /sn:0 {0}(1021,306)(1021,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w26;    //: /sn:0 {0}(368,306)(368,321){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w143;    //: /sn:0 {0}(910,306)(910,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w278;    //: /sn:0 {0}(1652,306)(1652,321){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w159;    //: /sn:0 {0}(1007,306)(1007,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w141;    //: /sn:0 {0}(917,306)(917,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w10;    //: /sn:0 {0}(254,214)(988,214)(988,290)(1003,290){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(935,156){13}
//: {14}(#:939,156)(1025,156){15}
//: {16}(#:1029,156)(1118,156){17}
//: {18}(#:1122,156)(1208,156){19}
//: {20}(#:1212,156)(1297,156){21}
//: {22}(#:1301,156)(1391,156){23}
//: {24}(#:1395,156)(1481,156){25}
//: {26}(#:1485,156)(1564,156){27}
//: {28}(#:1568,156)(1645,156){29}
//: {30}(#:1649,156)(1726,156)(1726,277){31}
//: {32}(1647,158)(1647,277){33}
//: {34}(1566,158)(1566,277){35}
//: {36}(1483,158)(1483,277){37}
//: {38}(1393,158)(1393,277){39}
//: {40}(1299,158)(1299,277){41}
//: {42}(1210,158)(1210,277){43}
//: {44}(1120,158)(1120,277){45}
//: {46}(1027,158)(1027,277){47}
//: {48}(937,158)(937,277){49}
//: {50}(842,158)(842,277){51}
//: {52}(744,158)(744,277){53}
//: {54}(649,158)(649,277){55}
//: {56}(560,158)(560,277){57}
//: {58}(459,158)(459,277){59}
//: {60}(363,158)(363,277){61}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w290;    //: /sn:0 {0}(1752,306)(1752,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w80;    //: /sn:0 {0}(654,306)(654,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire w277;    //: /sn:0 {0}(1655,306)(1655,321){1}
wire w149;    //: /sn:0 {0}(1042,306)(1042,321){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w160;    //: /sn:0 {0}(1004,306)(1004,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire w133;    //: /sn:0 {0}(945,306)(945,321){1}
wire w77;    //: /sn:0 {0}(664,306)(664,321){1}
wire w51;    //: /sn:0 {0}(439,306)(439,321){1}
//: enddecls

  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 53 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(w26), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(w33), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 61 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 37 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 50 ]
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(w269));   //: @(1566,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w1) @(1210, 156) /w:[ 20 -1 19 42 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 56 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 54 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g29 (w1) @(1120, 156) /w:[ 18 -1 17 44 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 52 ]
  _GGDECODER16 #(6, 6) g10 (.I(w1), .E(w11), .Z0(w128), .Z1(w129), .Z2(w130), .Z3(w131), .Z4(w132), .Z5(w133), .Z6(w134), .Z7(w135), .Z8(w136), .Z9(w137), .Z10(w138), .Z11(w139), .Z12(w140), .Z13(w141), .Z14(w142), .Z15(w143));   //: @(937,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(w69), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 57 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 30 -1 29 32 ]
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 51 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(w77), .Z4(w78), .Z5(w79), .Z6(w80), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(w85), .Z12(w86), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 55 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w1) @(1299, 156) /w:[ 22 -1 21 40 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 58 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: joint g33 (w1) @(1483, 156) /w:[ 26 -1 25 36 ]
  _GGDECODER16 #(6, 6) g12 (.I(w1), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g34 (w1) @(1566, 156) /w:[ 28 -1 27 34 ]
  //: joint g28 (w1) @(1027, 156) /w:[ 16 -1 15 46 ]
  _GGDECODER16 #(6, 6) g14 (.I(w1), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g11 (.I(w1), .E(w10), .Z0(w146), .Z1(w147), .Z2(w148), .Z3(w149), .Z4(w150), .Z5(w151), .Z6(w152), .Z7(w153), .Z8(w154), .Z9(w155), .Z10(w156), .Z11(w157), .Z12(w158), .Z13(w159), .Z14(w160), .Z15(w161));   //: @(1027,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(w44), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(w51), .Z14(w52), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 59 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 60 ]
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(w290), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 31 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g32 (w1) @(1393, 156) /w:[ 24 -1 23 38 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w1), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: joint g27 (w1) @(937, 156) /w:[ 14 -1 13 48 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w1), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 43 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin flags
module flags(x0_carry_flag, x2_parity_Overflow_flag, x7_sign_flag, x7_change_sign_flag, Flag_output, x1_change_Subtract_flag, x1_subtract_flag, x2_change_Parity_Overflow_flag, x4_change_Half_carry_flag, x0_change_carry_flag, x6_zero_flag, Flag_input, x6_change_zero_flag, x4_half_carry_flag);
//: interface  /sz:(405, 236) /bd:[ Li0>x7_sign_flag(192/236) Li1>x7_change_sign_flag(176/236) Li2>x6_zero_flag(160/236) Li3>x6_change_zero_flag(144/236) Li4>x4_half_carry_flag(128/236) Li5>x4_change_Half_carry_flag(112/236) Li6>x2_change_Parity_Overflow_flag(96/236) Li7>x2_parity_Overflow_flag(80/236) Li8>x1_subtract_flag(64/236) Li9>x1_change_Subtract_flag(48/236) Li10>x0_change_carry_flag(32/236) Li11>x0_carry_flag(16/236) Bi0>Flag_input[7:0](255/405) Bo0<Flag_output[7:0](110/405) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input x1_subtract_flag;    //: /sn:0 {0}(-10,-51)(128,-51){1}
input x0_carry_flag;    //: /sn:0 {0}(-10,-159)(52,-159)(52,-147){1}
input x4_half_carry_flag;    //: /sn:0 {0}(-10,242)(365,242){1}
input x7_sign_flag;    //: /sn:0 {0}(-11,460)(455,460)(455,473){1}
input x6_zero_flag;    //: /sn:0 {0}(407,362)(407,324)(-10,324){1}
input [7:0] Flag_input;    //: /sn:0 {0}(#:313,-191)(313,-240)(313,-240)(#:313,-291){1}
input x7_change_sign_flag;    //: /sn:0 {0}(-11,489)(442,489){1}
output [7:0] Flag_output;    //: /sn:0 {0}(#:313,572)(313,609)(313,609)(313,649){1}
input x1_change_Subtract_flag;    //: /sn:0 {0}(-10,-79)(141,-79)(141,-67){1}
input x4_change_Half_carry_flag;    //: /sn:0 {0}(378,226)(378,214)(-10,214){1}
input x2_change_Parity_Overflow_flag;    //: /sn:0 {0}(-10,70)(233,70){1}
input x2_parity_Overflow_flag;    //: /sn:0 {0}(-10,42)(246,42)(246,54){1}
input x0_change_carry_flag;    //: /sn:0 {0}(-10,-131)(39,-131){1}
input x6_change_zero_flag;    //: /sn:0 {0}(-10,378)(394,378){1}
wire w6;    //: /sn:0 {0}(328,566)(328,-185){1}
wire w7;    //: /sn:0 {0}(417,391)(417,400)(338,400)(338,566){1}
wire w4;    //: /sn:0 {0}(308,-185)(308,566){1}
wire w0;    //: /sn:0 {0}(62,-118)(62,162)(278,162)(278,566){1}
wire w3;    //: /sn:0 {0}(256,83)(256,139)(298,139)(298,566){1}
wire w22;    //: /sn:0 {0}(318,566)(318,270)(388,270)(388,255){1}
wire w19;    //: /sn:0 {0}(266,54)(266,-70)(298,-70)(298,-185){1}
wire w23;    //: /sn:0 {0}(427,362)(427,-57)(338,-57)(338,-185){1}
wire w24;    //: /sn:0 {0}(475,473)(475,-84)(348,-84)(348,-185){1}
wire w1;    //: /sn:0 {0}(151,-38)(151,152)(288,152)(288,566){1}
wire w8;    //: /sn:0 {0}(398,226)(398,160)(318,160)(318,-185){1}
wire w17;    //: /sn:0 {0}(161,-67)(161,-136)(288,-136)(288,-185){1}
wire w2;    //: /sn:0 {0}(72,-147)(72,-170)(278,-170)(278,-185){1}
wire w5;    //: /sn:0 {0}(348,566)(348,517)(465,517)(465,502){1}
//: enddecls

  //: IN g4 (x0_carry_flag) @(-12,-159) /sn:0 /w:[ 0 ]
  //: IN g8 (x2_parity_Overflow_flag) @(-12,42) /sn:0 /w:[ 0 ]
  _GGMUX2 #(8, 8) g3 (.I0(w8), .I1(x4_change_Half_carry_flag), .S(x4_half_carry_flag), .Z(w22));   //: @(388,242) /sn:0 /w:[ 0 0 1 1 ] /ss:0 /do:1
  //: IN g16 (x7_sign_flag) @(-13,460) /sn:0 /w:[ 0 ]
  //: IN g17 (x7_change_sign_flag) @(-13,489) /sn:0 /w:[ 0 ]
  //: OUT g2 (Flag_output) @(313,646) /sn:0 /R:3 /w:[ 1 ]
  _GGMUX2 #(8, 8) g1 (.I0(w17), .I1(x1_change_Subtract_flag), .S(x1_subtract_flag), .Z(w1));   //: @(151,-51) /sn:0 /w:[ 0 1 1 0 ] /ss:0 /do:1
  assign {w24, w23, w6, w8, w4, w19, w17, w2} = Flag_input; //: CONCAT g18  @(313,-190) /sn:0 /R:1 /w:[ 1 1 1 1 0 1 1 1 0 ] /dr:1 /tp:0 /drp:0
  assign Flag_output = {w5, w7, w6, w22, w4, w3, w1, w0}; //: CONCAT g10  @(313,571) /sn:0 /R:3 /w:[ 0 0 1 0 0 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: IN g6 (x1_change_Subtract_flag) @(-12,-79) /sn:0 /w:[ 0 ]
  //: IN g7 (x1_subtract_flag) @(-12,-51) /sn:0 /w:[ 0 ]
  //: IN g9 (x2_change_Parity_Overflow_flag) @(-12,70) /sn:0 /w:[ 0 ]
  _GGMUX2 #(8, 8) g22 (.I0(w2), .I1(x0_carry_flag), .S(x0_change_carry_flag), .Z(w0));   //: @(62,-131) /sn:0 /w:[ 0 1 1 0 ] /ss:0 /do:1
  _GGMUX2 #(8, 8) g33 (.I0(w23), .I1(x6_zero_flag), .S(x6_change_zero_flag), .Z(w7));   //: @(417,378) /sn:0 /w:[ 0 0 1 0 ] /ss:0 /do:1
  //: IN g12 (x4_change_Half_carry_flag) @(-12,214) /sn:0 /w:[ 1 ]
  _GGMUX2 #(8, 8) g28 (.I0(w19), .I1(x2_parity_Overflow_flag), .S(x2_change_Parity_Overflow_flag), .Z(w3));   //: @(256,70) /sn:0 /w:[ 0 1 1 0 ] /ss:0 /do:1
  _GGMUX2 #(8, 8) g34 (.I0(w24), .I1(x7_sign_flag), .S(x7_change_sign_flag), .Z(w5));   //: @(465,489) /sn:0 /w:[ 0 1 1 1 ] /ss:0 /do:1
  //: IN g5 (x0_change_carry_flag) @(-12,-131) /sn:0 /w:[ 0 ]
  //: IN g14 (x6_zero_flag) @(-12,324) /sn:0 /w:[ 1 ]
  //: IN g0 (Flag_input) @(313,-293) /sn:0 /R:3 /w:[ 1 ]
  //: IN g15 (x6_change_zero_flag) @(-12,378) /sn:0 /w:[ 0 ]
  //: IN g13 (x4_half_carry_flag) @(-12,242) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin instruction_IY_BITS
module instruction_IY_BITS(Instruction_input);
//: interface  /sz:(333, 534) /bd:[ Li0>Instruction_input[7:0](213/534) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w58;    //: /sn:0 {0}(579,306)(579,321){1}
wire w139;    //: /sn:0 {0}(924,306)(924,321){1}
wire w248;    //: /sn:0 {0}(1467,306)(1467,321){1}
wire w240;    //: /sn:0 {0}(1495,306)(1495,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w4;    //: /sn:0 {0}(254,193)(1527,193)(1527,290)(1542,290){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w282;    //: /sn:0 {0}(1638,306)(1638,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w303;    //: /sn:0 {0}(1706,306)(1706,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire w128;    //: /sn:0 {0}(963,306)(963,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w261;    //: /sn:0 {0}(1567,306)(1567,321){1}
wire w20;    //: /sn:0 {0}(389,306)(389,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w42;    //: /sn:0 {0}(471,306)(471,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w86;    //: /sn:0 {0}(633,306)(633,321){1}
wire w247;    //: /sn:0 {0}(1470,306)(1470,321){1}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w250;    //: /sn:0 {0}(1460,306)(1460,321){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w68;    //: /sn:0 {0}(544,306)(544,321){1}
wire w32;    //: /sn:0 {0}(347,306)(347,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w281;    //: /sn:0 {0}(1641,306)(1641,321){1}
wire w53;    //: /sn:0 {0}(432,306)(432,321){1}
wire w140;    //: /sn:0 {0}(921,306)(921,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w147;    //: /sn:0 {0}(1049,306)(1049,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w89;    //: /sn:0 {0}(622,306)(622,321){1}
wire w276;    //: /sn:0 {0}(1659,306)(1659,321){1}
wire w263;    //: /sn:0 {0}(1560,306)(1560,321){1}
wire w260;    //: /sn:0 {0}(1571,306)(1571,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w44;    //: /sn:0 {0}(464,306)(464,321){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w135;    //: /sn:0 {0}(938,306)(938,321){1}
wire w28;    //: /sn:0 {0}(361,306)(361,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w14;    //: /sn:0 {0}(254,228)(610,228)(610,290)(625,290){1}
wire w243;    //: /sn:0 {0}(1484,306)(1484,321){1}
wire w45;    //: /sn:0 {0}(460,306)(460,321){1}
wire w11;    //: /sn:0 {0}(254,218)(898,218)(898,290)(913,290){1}
wire w2;    //: /sn:0 {0}(254,186)(1687,186)(1687,290)(1702,290){1}
wire w74;    //: /sn:0 {0}(675,306)(675,321){1}
wire w78;    //: /sn:0 {0}(661,306)(661,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w296;    //: /sn:0 {0}(1731,306)(1731,321){1}
wire w129;    //: /sn:0 {0}(959,306)(959,321){1}
wire w274;    //: /sn:0 {0}(1666,306)(1666,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w15;    //: /sn:0 {0}(254,232)(521,232)(521,290)(536,290){1}
wire w272;    //: /sn:0 {0}(1673,306)(1673,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w87;    //: /sn:0 {0}(629,306)(629,321){1}
wire w43;    //: /sn:0 {0}(467,306)(467,321){1}
wire w286;    //: /sn:0 {0}(1624,306)(1624,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w40;    //: /sn:0 {0}(478,306)(478,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w262;    //: /sn:0 {0}(1564,306)(1564,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w264;    //: /sn:0 {0}(1557,306)(1557,321){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w34;    //: /sn:0 {0}(340,306)(340,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w158;    //: /sn:0 {0}(1011,306)(1011,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w62;    //: /sn:0 {0}(565,306)(565,321){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w241;    //: /sn:0 {0}(1491,306)(1491,321){1}
wire w142;    //: /sn:0 {0}(914,306)(914,321){1}
wire w299;    //: /sn:0 {0}(1720,306)(1720,321){1}
wire w82;    //: /sn:0 {0}(647,306)(647,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w148;    //: /sn:0 {0}(1046,306)(1046,321){1}
wire w71;    //: /sn:0 {0}(533,306)(533,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w154;    //: /sn:0 {0}(1025,306)(1025,321){1}
wire w156;    //: /sn:0 {0}(1018,306)(1018,321){1}
wire w255;    //: /sn:0 {0}(1588,306)(1588,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w66;    //: /sn:0 {0}(551,306)(551,321){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w63;    //: /sn:0 {0}(561,306)(561,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w130;    //: /sn:0 {0}(956,306)(956,321){1}
wire w285;    //: /sn:0 {0}(1627,306)(1627,321){1}
wire w21;    //: /sn:0 {0}(385,306)(385,321){1}
wire w256;    //: /sn:0 {0}(1585,306)(1585,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w131;    //: /sn:0 {0}(952,306)(952,321){1}
wire w268;    //: /sn:0 {0}(1543,306)(1543,321){1}
wire w246;    //: /sn:0 {0}(1474,306)(1474,321){1}
wire w293;    //: /sn:0 {0}(1741,306)(1741,321){1}
wire w302;    //: /sn:0 {0}(1710,306)(1710,321){1}
wire w304;    //: /sn:0 {0}(1703,306)(1703,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w52;    //: /sn:0 {0}(436,306)(436,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w244;    //: /sn:0 {0}(1481,306)(1481,321){1}
wire w75;    //: /sn:0 {0}(671,306)(671,321){1}
wire w150;    //: /sn:0 {0}(1039,306)(1039,321){1}
wire w33;    //: /sn:0 {0}(343,306)(343,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w69;    //: /sn:0 {0}(540,306)(540,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w300;    //: /sn:0 {0}(1717,306)(1717,321){1}
wire w257;    //: /sn:0 {0}(1581,306)(1581,321){1}
wire w47;    //: /sn:0 {0}(453,306)(453,321){1}
wire w146;    //: /sn:0 {0}(1053,306)(1053,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w294;    //: /sn:0 {0}(1738,306)(1738,321){1}
wire w245;    //: /sn:0 {0}(1477,306)(1477,321){1}
wire w85;    //: /sn:0 {0}(636,306)(636,321){1}
wire w151;    //: /sn:0 {0}(1035,306)(1035,321){1}
wire w161;    //: /sn:0 {0}(1000,306)(1000,321){1}
wire w297;    //: /sn:0 {0}(1727,306)(1727,321){1}
wire w137;    //: /sn:0 {0}(931,306)(931,321){1}
wire w267;    //: /sn:0 {0}(1546,306)(1546,321){1}
wire w238;    //: /sn:0 {0}(1502,306)(1502,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w38;    //: /sn:0 {0}(485,306)(485,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w265;    //: /sn:0 {0}(1553,306)(1553,321){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
wire w79;    //: /sn:0 {0}(657,306)(657,321){1}
wire w157;    //: /sn:0 {0}(1014,306)(1014,321){1}
wire w292;    //: /sn:0 {0}(1745,306)(1745,321){1}
wire w16;    //: /sn:0 {0}(254,235)(420,235)(420,290)(435,290){1}
wire w249;    //: /sn:0 {0}(1463,306)(1463,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w275;    //: /sn:0 {0}(1662,306)(1662,321){1}
wire w242;    //: /sn:0 {0}(1488,306)(1488,321){1}
wire w295;    //: /sn:0 {0}(1734,306)(1734,321){1}
wire w236;    //: /sn:0 {0}(1509,306)(1509,321){1}
wire w88;    //: /sn:0 {0}(626,306)(626,321){1}
wire w50;    //: /sn:0 {0}(443,306)(443,321){1}
wire w259;    //: /sn:0 {0}(1574,306)(1574,321){1}
wire w81;    //: /sn:0 {0}(650,306)(650,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w39;    //: /sn:0 {0}(481,306)(481,321){1}
wire w56;    //: /sn:0 {0}(586,306)(586,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w237;    //: /sn:0 {0}(1505,306)(1505,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w132;    //: /sn:0 {0}(949,306)(949,321){1}
wire w3;    //: /sn:0 {0}(254,190)(1608,190)(1608,290)(1623,290){1}
wire w22;    //: /sn:0 {0}(382,306)(382,321){1}
wire w273;    //: /sn:0 {0}(1669,306)(1669,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w30;    //: /sn:0 {0}(354,306)(354,321){1}
wire w29;    //: /sn:0 {0}(357,306)(357,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w152;    //: /sn:0 {0}(1032,306)(1032,321){1}
wire w138;    //: /sn:0 {0}(928,306)(928,321){1}
wire w269;    //: /sn:0 {0}(1539,306)(1539,321){1}
wire w31;    //: /sn:0 {0}(350,306)(350,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w266;    //: /sn:0 {0}(1550,306)(1550,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w46;    //: /sn:0 {0}(457,306)(457,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w67;    //: /sn:0 {0}(547,306)(547,321){1}
wire w136;    //: /sn:0 {0}(935,306)(935,321){1}
wire w134;    //: /sn:0 {0}(942,306)(942,321){1}
wire w35;    //: /sn:0 {0}(336,306)(336,321){1}
wire w284;    //: /sn:0 {0}(1631,306)(1631,321){1}
wire w41;    //: /sn:0 {0}(474,306)(474,321){1}
wire w153;    //: /sn:0 {0}(1028,306)(1028,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w283;    //: /sn:0 {0}(1634,306)(1634,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w155;    //: /sn:0 {0}(1021,306)(1021,321){1}
wire w305;    //: /sn:0 {0}(1699,306)(1699,321){1}
wire w83;    //: /sn:0 {0}(643,306)(643,321){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w254;    //: /sn:0 {0}(1592,306)(1592,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w26;    //: /sn:0 {0}(368,306)(368,321){1}
wire w76;    //: /sn:0 {0}(668,306)(668,321){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w279;    //: /sn:0 {0}(1648,306)(1648,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w65;    //: /sn:0 {0}(554,306)(554,321){1}
wire w143;    //: /sn:0 {0}(910,306)(910,321){1}
wire w251;    //: /sn:0 {0}(1456,306)(1456,321){1}
wire w291;    //: /sn:0 {0}(1748,306)(1748,321){1}
wire w59;    //: /sn:0 {0}(575,306)(575,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w278;    //: /sn:0 {0}(1652,306)(1652,321){1}
wire w239;    //: /sn:0 {0}(1498,306)(1498,321){1}
wire w25;    //: /sn:0 {0}(371,306)(371,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w159;    //: /sn:0 {0}(1007,306)(1007,321){1}
wire w60;    //: /sn:0 {0}(572,306)(572,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w141;    //: /sn:0 {0}(917,306)(917,321){1}
wire w258;    //: /sn:0 {0}(1578,306)(1578,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w10;    //: /sn:0 {0}(254,214)(988,214)(988,290)(1003,290){1}
wire w23;    //: /sn:0 {0}(378,306)(378,321){1}
wire w70;    //: /sn:0 {0}(537,306)(537,321){1}
wire w84;    //: /sn:0 {0}(640,306)(640,321){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w24;    //: /sn:0 {0}(375,306)(375,321){1}
wire [3:0] w1;    //: /sn:0 {0}(#:363,128)(363,154){1}
//: {2}(#:365,156)(457,156){3}
//: {4}(#:461,156)(558,156){5}
//: {6}(#:562,156)(647,156){7}
//: {8}(#:651,156)(742,156){9}
//: {10}(#:746,156)(840,156){11}
//: {12}(#:844,156)(935,156){13}
//: {14}(#:939,156)(1025,156){15}
//: {16}(#:1029,156)(1118,156){17}
//: {18}(#:1122,156)(1208,156){19}
//: {20}(#:1212,156)(1297,156){21}
//: {22}(#:1301,156)(1391,156){23}
//: {24}(#:1395,156)(1481,156){25}
//: {26}(#:1485,156)(1564,156){27}
//: {28}(#:1568,156)(1645,156){29}
//: {30}(#:1649,156)(1726,156)(1726,277){31}
//: {32}(1647,158)(1647,277){33}
//: {34}(1566,158)(1566,277){35}
//: {36}(1483,158)(1483,277){37}
//: {38}(1393,158)(1393,277){39}
//: {40}(1299,158)(1299,277){41}
//: {42}(1210,158)(1210,277){43}
//: {44}(1120,158)(1120,277){45}
//: {46}(1027,158)(1027,277){47}
//: {48}(937,158)(937,277){49}
//: {50}(842,158)(842,277){51}
//: {52}(744,158)(744,277){53}
//: {54}(649,158)(649,277){55}
//: {56}(560,158)(560,277){57}
//: {58}(459,158)(459,277){59}
//: {60}(363,158)(363,277){61}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w287;    //: /sn:0 {0}(1620,306)(1620,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w290;    //: /sn:0 {0}(1752,306)(1752,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w27;    //: /sn:0 {0}(364,306)(364,321){1}
wire w17;    //: /sn:0 {0}(254,239)(324,239)(324,290)(339,290){1}
wire w80;    //: /sn:0 {0}(654,306)(654,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w49;    //: /sn:0 {0}(446,306)(446,321){1}
wire w48;    //: /sn:0 {0}(450,306)(450,321){1}
wire w280;    //: /sn:0 {0}(1645,306)(1645,321){1}
wire w277;    //: /sn:0 {0}(1655,306)(1655,321){1}
wire w149;    //: /sn:0 {0}(1042,306)(1042,321){1}
wire w61;    //: /sn:0 {0}(568,306)(568,321){1}
wire w5;    //: /sn:0 {0}(254,197)(1444,197)(1444,290)(1459,290){1}
wire w64;    //: /sn:0 {0}(558,306)(558,321){1}
wire w160;    //: /sn:0 {0}(1004,306)(1004,321){1}
wire w298;    //: /sn:0 {0}(1724,306)(1724,321){1}
wire w301;    //: /sn:0 {0}(1713,306)(1713,321){1}
wire w57;    //: /sn:0 {0}(582,306)(582,321){1}
wire w133;    //: /sn:0 {0}(945,306)(945,321){1}
wire w77;    //: /sn:0 {0}(664,306)(664,321){1}
wire w51;    //: /sn:0 {0}(439,306)(439,321){1}
//: enddecls

  _GGDECODER16 #(6, 6) g8 (.I(w1), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 53 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g4 (.I(w1), .E(w17), .Z0(w20), .Z1(w21), .Z2(w22), .Z3(w23), .Z4(w24), .Z5(w25), .Z6(w26), .Z7(w27), .Z8(w28), .Z9(w29), .Z10(w30), .Z11(w31), .Z12(w32), .Z13(w33), .Z14(w34), .Z15(w35));   //: @(363,290) /sn:0 /w:[ 61 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g16 (.I(w1), .E(w5), .Z0(w236), .Z1(w237), .Z2(w238), .Z3(w239), .Z4(w240), .Z5(w241), .Z6(w242), .Z7(w243), .Z8(w244), .Z9(w245), .Z10(w246), .Z11(w247), .Z12(w248), .Z13(w249), .Z14(w250), .Z15(w251));   //: @(1483,290) /sn:0 /w:[ 37 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(842, 156) /w:[ 12 -1 11 50 ]
  _GGDECODER16 #(6, 6) g17 (.I(w1), .E(w4), .Z0(w254), .Z1(w255), .Z2(w256), .Z3(w257), .Z4(w258), .Z5(w259), .Z6(w260), .Z7(w261), .Z8(w262), .Z9(w263), .Z10(w264), .Z11(w265), .Z12(w266), .Z13(w267), .Z14(w268), .Z15(w269));   //: @(1566,290) /sn:0 /w:[ 35 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w1) @(1210, 156) /w:[ 20 -1 19 42 ]
  //: joint g23 (w1) @(560, 156) /w:[ 6 -1 5 56 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  //: joint g24 (w1) @(649, 156) /w:[ 8 -1 7 54 ]
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g29 (w1) @(1120, 156) /w:[ 18 -1 17 44 ]
  _GGDECODER16 #(6, 6) g18 (.I(w1), .E(w3), .Z0(w272), .Z1(w273), .Z2(w274), .Z3(w275), .Z4(w276), .Z5(w277), .Z6(w278), .Z7(w279), .Z8(w280), .Z9(w281), .Z10(w282), .Z11(w283), .Z12(w284), .Z13(w285), .Z14(w286), .Z15(w287));   //: @(1647,290) /sn:0 /w:[ 33 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g25 (w1) @(744, 156) /w:[ 10 -1 9 52 ]
  _GGDECODER16 #(6, 6) g10 (.I(w1), .E(w11), .Z0(w128), .Z1(w129), .Z2(w130), .Z3(w131), .Z4(w132), .Z5(w133), .Z6(w134), .Z7(w135), .Z8(w136), .Z9(w137), .Z10(w138), .Z11(w139), .Z12(w140), .Z13(w141), .Z14(w142), .Z15(w143));   //: @(937,290) /sn:0 /w:[ 49 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g6 (.I(w1), .E(w15), .Z0(w56), .Z1(w57), .Z2(w58), .Z3(w59), .Z4(w60), .Z5(w61), .Z6(w62), .Z7(w63), .Z8(w64), .Z9(w65), .Z10(w66), .Z11(w67), .Z12(w68), .Z13(w69), .Z14(w70), .Z15(w71));   //: @(560,290) /sn:0 /w:[ 57 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g35 (w1) @(1647, 156) /w:[ 30 -1 29 32 ]
  _GGDECODER16 #(6, 6) g9 (.I(w1), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 51 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g7 (.I(w1), .E(w14), .Z0(w74), .Z1(w75), .Z2(w76), .Z3(w77), .Z4(w78), .Z5(w79), .Z6(w80), .Z7(w81), .Z8(w82), .Z9(w83), .Z10(w84), .Z11(w85), .Z12(w86), .Z13(w87), .Z14(w88), .Z15(w89));   //: @(649,290) /sn:0 /w:[ 55 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w1) @(1299, 156) /w:[ 22 -1 21 40 ]
  //: joint g22 (w1) @(459, 156) /w:[ 4 -1 3 58 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  //: joint g33 (w1) @(1483, 156) /w:[ 26 -1 25 36 ]
  _GGDECODER16 #(6, 6) g12 (.I(w1), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 45 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g34 (w1) @(1566, 156) /w:[ 28 -1 27 34 ]
  //: joint g28 (w1) @(1027, 156) /w:[ 16 -1 15 46 ]
  _GGDECODER16 #(6, 6) g14 (.I(w1), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 41 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g11 (.I(w1), .E(w10), .Z0(w146), .Z1(w147), .Z2(w148), .Z3(w149), .Z4(w150), .Z5(w151), .Z6(w152), .Z7(w153), .Z8(w154), .Z9(w155), .Z10(w156), .Z11(w157), .Z12(w158), .Z13(w159), .Z14(w160), .Z15(w161));   //: @(1027,290) /sn:0 /w:[ 47 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  _GGDECODER16 #(6, 6) g5 (.I(w1), .E(w16), .Z0(w38), .Z1(w39), .Z2(w40), .Z3(w41), .Z4(w42), .Z5(w43), .Z6(w44), .Z7(w45), .Z8(w46), .Z9(w47), .Z10(w48), .Z11(w49), .Z12(w50), .Z13(w51), .Z14(w52), .Z15(w53));   //: @(459,290) /sn:0 /w:[ 59 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g21 (w1) @(363, 156) /w:[ 2 1 -1 60 ]
  _GGDECODER16 #(6, 6) g19 (.I(w1), .E(w2), .Z0(w290), .Z1(w291), .Z2(w292), .Z3(w293), .Z4(w294), .Z5(w295), .Z6(w296), .Z7(w297), .Z8(w298), .Z9(w299), .Z10(w300), .Z11(w301), .Z12(w302), .Z13(w303), .Z14(w304), .Z15(w305));   //: @(1726,290) /sn:0 /w:[ 31 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g32 (w1) @(1393, 156) /w:[ 24 -1 23 38 ]
  assign w1 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w1), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 39 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: joint g27 (w1) @(937, 156) /w:[ 14 -1 13 48 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w1), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 43 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

//: /netlistBegin instruction_EXTD
module instruction_EXTD(Instruction_input);
//: interface  /sz:(315, 456) /bd:[ Li0>Instruction_input[7:0](182/456) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w18;    //: /sn:0 {0}(168,204)(168,250)(238,250)(238,235){1}
input [7:0] Instruction_input;    //: /sn:0 {0}(#:170,124)(197,124){1}
//: {2}(198,124)(362,124){3}
//: {4}(363,124)(413,124){5}
wire w207;    //: /sn:0 {0}(1300,306)(1300,321){1}
wire w6;    //: /sn:0 {0}(254,200)(1354,200)(1354,290)(1369,290){1}
wire w16;    //: /sn:0 {0}(254,235)(415,235)(415,384){1}
wire w183;    //: /sn:0 {0}(1232,306)(1232,321){1}
wire w13;    //: /sn:0 {0}(254,225)(705,225)(705,290)(720,290){1}
wire w114;    //: /sn:0 {0}(854,306)(854,321){1}
wire w7;    //: /sn:0 {0}(254,204)(1260,204)(1260,290)(1275,290){1}
wire w174;    //: /sn:0 {0}(1111,306)(1111,321){1}
wire w192;    //: /sn:0 {0}(1201,306)(1201,321){1}
wire w197;    //: /sn:0 {0}(1183,306)(1183,321){1}
wire w171;    //: /sn:0 {0}(1121,306)(1121,321){1}
wire w205;    //: /sn:0 {0}(1307,306)(1307,321){1}
wire w165;    //: /sn:0 {0}(1142,306)(1142,321){1}
wire w203;    //: /sn:0 {0}(1314,306)(1314,321){1}
wire w175;    //: /sn:0 {0}(1107,306)(1107,321){1}
wire w229;    //: /sn:0 {0}(1380,306)(1380,321){1}
wire w25;    //: /sn:0 {0}(254,228)(425,228)(425,384){1}
wire w186;    //: /sn:0 {0}(1222,306)(1222,321){1}
wire w123;    //: /sn:0 {0}(822,306)(822,321){1}
wire w177;    //: /sn:0 {0}(1100,306)(1100,321){1}
wire w202;    //: /sn:0 {0}(1318,306)(1318,321){1}
wire w101;    //: /sn:0 {0}(738,306)(738,321){1}
wire w164;    //: /sn:0 {0}(1146,306)(1146,321){1}
wire w223;    //: /sn:0 {0}(1401,306)(1401,321){1}
wire w117;    //: /sn:0 {0}(843,306)(843,321){1}
wire w176;    //: /sn:0 {0}(1104,306)(1104,321){1}
wire w189;    //: /sn:0 {0}(1211,306)(1211,321){1}
wire [3:0] w0;    //: /sn:0 {0}(#:198,128)(198,213)(225,213){1}
wire w22;    //: /sn:0 {0}(254,197)(440,197)(440,384){1}
wire w20;    //: /sn:0 {0}(433,434)(433,405){1}
wire w188;    //: /sn:0 {0}(1215,306)(1215,321){1}
wire w222;    //: /sn:0 {0}(1405,306)(1405,321){1}
wire w226;    //: /sn:0 {0}(1391,306)(1391,321){1}
wire w124;    //: /sn:0 {0}(819,306)(819,321){1}
wire w209;    //: /sn:0 {0}(1293,306)(1293,321){1}
wire w225;    //: /sn:0 {0}(1394,306)(1394,321){1}
wire w196;    //: /sn:0 {0}(1187,306)(1187,321){1}
wire w195;    //: /sn:0 {0}(1190,306)(1190,321){1}
wire w185;    //: /sn:0 {0}(1225,306)(1225,321){1}
wire w112;    //: /sn:0 {0}(861,306)(861,321){1}
wire w119;    //: /sn:0 {0}(836,306)(836,321){1}
wire w122;    //: /sn:0 {0}(826,306)(826,321){1}
wire w218;    //: /sn:0 {0}(1419,306)(1419,321){1}
wire w170;    //: /sn:0 {0}(1125,306)(1125,321){1}
wire w210;    //: /sn:0 {0}(1290,306)(1290,321){1}
wire w227;    //: /sn:0 {0}(1387,306)(1387,321){1}
wire w19;    //: /sn:0 {0}(254,190)(450,190)(450,384){1}
wire w190;    //: /sn:0 {0}(1208,306)(1208,321){1}
wire w12;    //: /sn:0 {0}(254,221)(803,221)(803,290)(818,290){1}
wire w168;    //: /sn:0 {0}(1132,306)(1132,321){1}
wire w214;    //: /sn:0 {0}(1276,306)(1276,321){1}
wire w206;    //: /sn:0 {0}(1304,306)(1304,321){1}
wire w178;    //: /sn:0 {0}(1097,306)(1097,321){1}
wire w211;    //: /sn:0 {0}(1286,306)(1286,321){1}
wire w23;    //: /sn:0 {0}(254,214)(435,214)(435,384){1}
wire w111;    //: /sn:0 {0}(864,306)(864,321){1}
wire w179;    //: /sn:0 {0}(1093,306)(1093,321){1}
wire w21;    //: /sn:0 {0}(254,193)(445,193)(445,384){1}
wire w24;    //: /sn:0 {0}(254,218)(430,218)(430,384){1}
wire [3:0] w108;    //: /sn:0 {0}(1393,277)(1393,156)(#:1301,156){1}
//: {2}(1297,156)(#:1212,156){3}
//: {4}(1208,156)(#:1122,156){5}
//: {6}(1118,156)(#:844,156){7}
//: {8}(840,156)(#:746,156){9}
//: {10}(742,156)(363,156)(#:363,128){11}
//: {12}(744,158)(744,277){13}
//: {14}(842,158)(842,277){15}
//: {16}(1120,158)(1120,277){17}
//: {18}(1210,158)(1210,277){19}
//: {20}(1299,158)(1299,277){21}
wire w106;    //: /sn:0 {0}(721,306)(721,321){1}
wire w121;    //: /sn:0 {0}(829,306)(829,321){1}
wire w201;    //: /sn:0 {0}(1321,306)(1321,321){1}
wire w1;    //: /sn:0 {0}(254,186)(455,186)(455,384){1}
wire w104;    //: /sn:0 {0}(728,306)(728,321){1}
wire w194;    //: /sn:0 {0}(1194,306)(1194,321){1}
wire w116;    //: /sn:0 {0}(847,306)(847,321){1}
wire w224;    //: /sn:0 {0}(1398,306)(1398,321){1}
wire w213;    //: /sn:0 {0}(1279,306)(1279,321){1}
wire w8;    //: /sn:0 {0}(254,207)(1171,207)(1171,290)(1186,290){1}
wire w115;    //: /sn:0 {0}(850,306)(850,321){1}
wire w230;    //: /sn:0 {0}(1377,306)(1377,321){1}
wire w110;    //: /sn:0 {0}(868,306)(868,321){1}
wire w182;    //: /sn:0 {0}(1236,306)(1236,321){1}
wire w200;    //: /sn:0 {0}(1325,306)(1325,321){1}
wire w95;    //: /sn:0 {0}(759,306)(759,321){1}
wire w232;    //: /sn:0 {0}(1370,306)(1370,321){1}
wire w233;    //: /sn:0 {0}(1366,306)(1366,321){1}
wire w191;    //: /sn:0 {0}(1204,306)(1204,321){1}
wire w103;    //: /sn:0 {0}(731,306)(731,321){1}
wire w98;    //: /sn:0 {0}(749,306)(749,321){1}
wire w167;    //: /sn:0 {0}(1135,306)(1135,321){1}
wire w193;    //: /sn:0 {0}(1197,306)(1197,321){1}
wire w17;    //: /sn:0 {0}(410,384)(410,239)(254,239){1}
wire w187;    //: /sn:0 {0}(1218,306)(1218,321){1}
wire w169;    //: /sn:0 {0}(1128,306)(1128,321){1}
wire w212;    //: /sn:0 {0}(1283,306)(1283,321){1}
wire w118;    //: /sn:0 {0}(840,306)(840,321){1}
wire w113;    //: /sn:0 {0}(857,306)(857,321){1}
wire w215;    //: /sn:0 {0}(1272,306)(1272,321){1}
wire w219;    //: /sn:0 {0}(1415,306)(1415,321){1}
wire w120;    //: /sn:0 {0}(833,306)(833,321){1}
wire w204;    //: /sn:0 {0}(1311,306)(1311,321){1}
wire w166;    //: /sn:0 {0}(1139,306)(1139,321){1}
wire w105;    //: /sn:0 {0}(724,306)(724,321){1}
wire w184;    //: /sn:0 {0}(1229,306)(1229,321){1}
wire w15;    //: /sn:0 {0}(254,232)(420,232)(420,384){1}
wire w228;    //: /sn:0 {0}(1384,306)(1384,321){1}
wire w94;    //: /sn:0 {0}(763,306)(763,321){1}
wire w92;    //: /sn:0 {0}(770,306)(770,321){1}
wire w102;    //: /sn:0 {0}(735,306)(735,321){1}
wire w173;    //: /sn:0 {0}(1114,306)(1114,321){1}
wire w172;    //: /sn:0 {0}(1118,306)(1118,321){1}
wire w231;    //: /sn:0 {0}(1373,306)(1373,321){1}
wire w9;    //: /sn:0 {0}(254,211)(1084,211)(1084,290)(1096,290){1}
wire w107;    //: /sn:0 {0}(717,306)(717,321){1}
wire w97;    //: /sn:0 {0}(752,306)(752,321){1}
wire w208;    //: /sn:0 {0}(1297,306)(1297,321){1}
wire w220;    //: /sn:0 {0}(1412,306)(1412,321){1}
wire w221;    //: /sn:0 {0}(1408,306)(1408,321){1}
wire w100;    //: /sn:0 {0}(742,306)(742,321){1}
wire w99;    //: /sn:0 {0}(745,306)(745,321){1}
wire w96;    //: /sn:0 {0}(756,306)(756,321){1}
wire w125;    //: /sn:0 {0}(815,306)(815,321){1}
wire w93;    //: /sn:0 {0}(766,306)(766,321){1}
//: enddecls

  _GGOR10 #(22) g4 (.I0(w1), .I1(w19), .I2(w21), .I3(w22), .I4(w23), .I5(w24), .I6(w25), .I7(w15), .I8(w16), .I9(w17), .Z(w20));   //: @(433,395) /sn:0 /R:3 /w:[ 1 1 1 1 1 1 1 1 1 0 1 ]
  _GGDECODER16 #(6, 6) g8 (.I(w108), .E(w13), .Z0(w92), .Z1(w93), .Z2(w94), .Z3(w95), .Z4(w96), .Z5(w97), .Z6(w98), .Z7(w99), .Z8(w100), .Z9(w101), .Z10(w102), .Z11(w103), .Z12(w104), .Z13(w105), .Z14(w106), .Z15(w107));   //: @(744,290) /sn:0 /w:[ 13 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: VDD g3 (w18) @(179,204) /sn:0 /w:[ 0 ]
  //: joint g26 (w108) @(842, 156) /w:[ 7 -1 8 14 ]
  assign w0 = Instruction_input[7:4]; //: TAP g2 @(198,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g30 (w108) @(1210, 156) /w:[ 3 -1 4 18 ]
  //: frame g39 @(1437,260) /sn:0 /wi:333 /ht:91 /tx:"0-63 (00-3F)"
  _GGDECODER16 #(6, 6) g1 (.I(w0), .E(w18), .Z0(w1), .Z1(w19), .Z2(w21), .Z3(w22), .Z4(w6), .Z5(w7), .Z6(w8), .Z7(w9), .Z8(w23), .Z9(w24), .Z10(w12), .Z11(w13), .Z12(w25), .Z13(w15), .Z14(w16), .Z15(w17));   //: @(238,213) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /ss:0 /do:1
  //: joint g29 (w108) @(1120, 156) /w:[ 5 -1 6 16 ]
  //: joint g25 (w108) @(744, 156) /w:[ 9 -1 10 12 ]
  _GGDECODER16 #(6, 6) g9 (.I(w108), .E(w12), .Z0(w110), .Z1(w111), .Z2(w112), .Z3(w113), .Z4(w114), .Z5(w115), .Z6(w116), .Z7(w117), .Z8(w118), .Z9(w119), .Z10(w120), .Z11(w121), .Z12(w122), .Z13(w123), .Z14(w124), .Z15(w125));   //: @(842,290) /sn:0 /w:[ 15 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: joint g31 (w108) @(1299, 156) /w:[ 1 -1 2 20 ]
  //: frame g36 @(300,259) /sn:0 /wi:388 /ht:92 /tx:"192-255 (C0-FF)"
  _GGDECODER16 #(6, 6) g12 (.I(w108), .E(w9), .Z0(w164), .Z1(w165), .Z2(w166), .Z3(w167), .Z4(w168), .Z5(w169), .Z6(w170), .Z7(w171), .Z8(w172), .Z9(w173), .Z10(w174), .Z11(w175), .Z12(w176), .Z13(w177), .Z14(w178), .Z15(w179));   //: @(1120,290) /sn:0 /w:[ 17 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: LED g5 (w20) @(433,441) /sn:0 /R:2 /w:[ 0 ] /type:0
  _GGDECODER16 #(6, 6) g14 (.I(w108), .E(w7), .Z0(w200), .Z1(w201), .Z2(w202), .Z3(w203), .Z4(w204), .Z5(w205), .Z6(w206), .Z7(w207), .Z8(w208), .Z9(w209), .Z10(w210), .Z11(w211), .Z12(w212), .Z13(w213), .Z14(w214), .Z15(w215));   //: @(1299,290) /sn:0 /w:[ 21 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  assign w108 = Instruction_input[3:0]; //: TAP g20 @(363,122) /sn:0 /R:1 /w:[ 11 3 4 ] /ss:1
  //: frame g38 @(1075,259) /sn:0 /wi:354 /ht:92 /tx:"64-127 (40-7F)"
  _GGDECODER16 #(6, 6) g15 (.I(w108), .E(w6), .Z0(w218), .Z1(w219), .Z2(w220), .Z3(w221), .Z4(w222), .Z5(w223), .Z6(w224), .Z7(w225), .Z8(w226), .Z9(w227), .Z10(w228), .Z11(w229), .Z12(w230), .Z13(w231), .Z14(w232), .Z15(w233));   //: @(1393,290) /sn:0 /w:[ 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1
  //: IN g0 (Instruction_input) @(168,124) /sn:0 /w:[ 0 ]
  //: frame g37 @(699,258) /sn:0 /wi:366 /ht:93 /tx:"128-191 (80-BF)"
  _GGDECODER16 #(6, 6) g13 (.I(w108), .E(w8), .Z0(w182), .Z1(w183), .Z2(w184), .Z3(w185), .Z4(w186), .Z5(w187), .Z6(w188), .Z7(w189), .Z8(w190), .Z9(w191), .Z10(w192), .Z11(w193), .Z12(w194), .Z13(w195), .Z14(w196), .Z15(w197));   //: @(1210,290) /sn:0 /w:[ 19 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /ss:0 /do:1

endmodule
//: /netlistEnd

